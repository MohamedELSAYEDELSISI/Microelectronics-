
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_Logix_control_rf is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_Logix_control_rf;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Logix_control_rf.all;

entity Logix_control_rf_DW01_incdec_1_DW01_incdec_2 is

   port( A : in std_logic_vector (31 downto 0);  INC_DEC : in std_logic;  SUM :
         out std_logic_vector (31 downto 0));

end Logix_control_rf_DW01_incdec_1_DW01_incdec_2;

architecture SYN_rpl of Logix_control_rf_DW01_incdec_1_DW01_incdec_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n2, n_1000, 
      n_1001 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => INC_DEC, CI => carry_31_port, CO =>
                           n_1000, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => INC_DEC, CI => carry_30_port, CO =>
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => INC_DEC, CI => carry_29_port, CO =>
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => INC_DEC, CI => carry_28_port, CO =>
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => INC_DEC, CI => carry_27_port, CO =>
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => INC_DEC, CI => carry_26_port, CO =>
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => INC_DEC, CI => carry_25_port, CO =>
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => INC_DEC, CI => carry_24_port, CO =>
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => INC_DEC, CI => carry_23_port, CO =>
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => INC_DEC, CI => carry_22_port, CO =>
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => INC_DEC, CI => carry_21_port, CO =>
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => INC_DEC, CI => carry_20_port, CO =>
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => INC_DEC, CI => carry_19_port, CO =>
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => INC_DEC, CI => carry_18_port, CO =>
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => INC_DEC, CI => carry_17_port, CO =>
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => INC_DEC, CI => carry_16_port, CO =>
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => INC_DEC, CI => carry_15_port, CO =>
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => INC_DEC, CI => carry_14_port, CO =>
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => INC_DEC, CI => carry_13_port, CO =>
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => INC_DEC, CI => carry_12_port, CO =>
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => INC_DEC, CI => carry_11_port, CO =>
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => INC_DEC, CI => carry_10_port, CO =>
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => INC_DEC, CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => INC_DEC, CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => INC_DEC, CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => INC_DEC, CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => INC_DEC, CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => INC_DEC, CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => INC_DEC, CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => INC_DEC, CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => INC_DEC, CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => INC_DEC, CI => n2, CO => carry_1_port
                           , S => n_1001);
   U1 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U2 : INV_X1 port map( A => INC_DEC, ZN => n2);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Logix_control_rf.all;

entity Logix_control_rf_DW01_incdec_0_DW01_incdec_1 is

   port( A : in std_logic_vector (31 downto 0);  INC_DEC : in std_logic;  SUM :
         out std_logic_vector (31 downto 0));

end Logix_control_rf_DW01_incdec_0_DW01_incdec_1;

architecture SYN_rpl of Logix_control_rf_DW01_incdec_0_DW01_incdec_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n2, n_1002, 
      n_1003 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => INC_DEC, CI => carry_31_port, CO =>
                           n_1002, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => INC_DEC, CI => carry_30_port, CO =>
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => INC_DEC, CI => carry_29_port, CO =>
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => INC_DEC, CI => carry_28_port, CO =>
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => INC_DEC, CI => carry_27_port, CO =>
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => INC_DEC, CI => carry_26_port, CO =>
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => INC_DEC, CI => carry_25_port, CO =>
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => INC_DEC, CI => carry_24_port, CO =>
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => INC_DEC, CI => carry_23_port, CO =>
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => INC_DEC, CI => carry_22_port, CO =>
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => INC_DEC, CI => carry_21_port, CO =>
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => INC_DEC, CI => carry_20_port, CO =>
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => INC_DEC, CI => carry_19_port, CO =>
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => INC_DEC, CI => carry_18_port, CO =>
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => INC_DEC, CI => carry_17_port, CO =>
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => INC_DEC, CI => carry_16_port, CO =>
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => INC_DEC, CI => carry_15_port, CO =>
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => INC_DEC, CI => carry_14_port, CO =>
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => INC_DEC, CI => carry_13_port, CO =>
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => INC_DEC, CI => carry_12_port, CO =>
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => INC_DEC, CI => carry_11_port, CO =>
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => INC_DEC, CI => carry_10_port, CO =>
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => INC_DEC, CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => INC_DEC, CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => INC_DEC, CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => INC_DEC, CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => INC_DEC, CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => INC_DEC, CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => INC_DEC, CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => INC_DEC, CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => INC_DEC, CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => INC_DEC, CI => n2, CO => carry_1_port
                           , S => n_1003);
   U1 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U2 : INV_X1 port map( A => INC_DEC, ZN => n2);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Logix_control_rf.all;

entity register_file_address_length5_Data_parallelism64 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_address_length5_Data_parallelism64;

architecture SYN_A of register_file_address_length5_Data_parallelism64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal REGISTERS_0_63_port, REGISTERS_0_62_port, REGISTERS_0_61_port, 
      REGISTERS_0_60_port, REGISTERS_0_59_port, REGISTERS_0_58_port, 
      REGISTERS_0_57_port, REGISTERS_0_56_port, REGISTERS_0_55_port, 
      REGISTERS_0_54_port, REGISTERS_0_53_port, REGISTERS_0_52_port, 
      REGISTERS_0_51_port, REGISTERS_0_50_port, REGISTERS_0_49_port, 
      REGISTERS_0_48_port, REGISTERS_0_47_port, REGISTERS_0_46_port, 
      REGISTERS_0_45_port, REGISTERS_0_44_port, REGISTERS_0_43_port, 
      REGISTERS_0_42_port, REGISTERS_0_41_port, REGISTERS_0_40_port, 
      REGISTERS_0_39_port, REGISTERS_0_38_port, REGISTERS_0_37_port, 
      REGISTERS_0_36_port, REGISTERS_0_35_port, REGISTERS_0_34_port, 
      REGISTERS_0_33_port, REGISTERS_0_32_port, REGISTERS_0_31_port, 
      REGISTERS_0_30_port, REGISTERS_0_29_port, REGISTERS_0_28_port, 
      REGISTERS_0_27_port, REGISTERS_0_26_port, REGISTERS_0_25_port, 
      REGISTERS_0_24_port, REGISTERS_0_23_port, REGISTERS_0_22_port, 
      REGISTERS_0_21_port, REGISTERS_0_20_port, REGISTERS_0_19_port, 
      REGISTERS_0_18_port, REGISTERS_0_17_port, REGISTERS_0_16_port, 
      REGISTERS_0_15_port, REGISTERS_0_14_port, REGISTERS_0_13_port, 
      REGISTERS_0_12_port, REGISTERS_0_11_port, REGISTERS_0_10_port, 
      REGISTERS_0_9_port, REGISTERS_0_8_port, REGISTERS_0_7_port, 
      REGISTERS_0_6_port, REGISTERS_0_5_port, REGISTERS_0_4_port, 
      REGISTERS_0_3_port, REGISTERS_0_2_port, REGISTERS_0_1_port, 
      REGISTERS_0_0_port, REGISTERS_1_63_port, REGISTERS_1_62_port, 
      REGISTERS_1_61_port, REGISTERS_1_60_port, REGISTERS_1_59_port, 
      REGISTERS_1_58_port, REGISTERS_1_57_port, REGISTERS_1_56_port, 
      REGISTERS_1_55_port, REGISTERS_1_54_port, REGISTERS_1_53_port, 
      REGISTERS_1_52_port, REGISTERS_1_51_port, REGISTERS_1_50_port, 
      REGISTERS_1_49_port, REGISTERS_1_48_port, REGISTERS_1_47_port, 
      REGISTERS_1_46_port, REGISTERS_1_45_port, REGISTERS_1_44_port, 
      REGISTERS_1_43_port, REGISTERS_1_42_port, REGISTERS_1_41_port, 
      REGISTERS_1_40_port, REGISTERS_1_39_port, REGISTERS_1_38_port, 
      REGISTERS_1_37_port, REGISTERS_1_36_port, REGISTERS_1_35_port, 
      REGISTERS_1_34_port, REGISTERS_1_33_port, REGISTERS_1_32_port, 
      REGISTERS_1_31_port, REGISTERS_1_30_port, REGISTERS_1_29_port, 
      REGISTERS_1_28_port, REGISTERS_1_27_port, REGISTERS_1_26_port, 
      REGISTERS_1_25_port, REGISTERS_1_24_port, REGISTERS_1_23_port, 
      REGISTERS_1_22_port, REGISTERS_1_21_port, REGISTERS_1_20_port, 
      REGISTERS_1_19_port, REGISTERS_1_18_port, REGISTERS_1_17_port, 
      REGISTERS_1_16_port, REGISTERS_1_15_port, REGISTERS_1_14_port, 
      REGISTERS_1_13_port, REGISTERS_1_12_port, REGISTERS_1_11_port, 
      REGISTERS_1_10_port, REGISTERS_1_9_port, REGISTERS_1_8_port, 
      REGISTERS_1_7_port, REGISTERS_1_6_port, REGISTERS_1_5_port, 
      REGISTERS_1_4_port, REGISTERS_1_3_port, REGISTERS_1_2_port, 
      REGISTERS_1_1_port, REGISTERS_1_0_port, REGISTERS_2_63_port, 
      REGISTERS_2_62_port, REGISTERS_2_61_port, REGISTERS_2_60_port, 
      REGISTERS_2_59_port, REGISTERS_2_58_port, REGISTERS_2_57_port, 
      REGISTERS_2_56_port, REGISTERS_2_55_port, REGISTERS_2_54_port, 
      REGISTERS_2_53_port, REGISTERS_2_52_port, REGISTERS_2_51_port, 
      REGISTERS_2_50_port, REGISTERS_2_49_port, REGISTERS_2_48_port, 
      REGISTERS_2_47_port, REGISTERS_2_46_port, REGISTERS_2_45_port, 
      REGISTERS_2_44_port, REGISTERS_2_43_port, REGISTERS_2_42_port, 
      REGISTERS_2_41_port, REGISTERS_2_40_port, REGISTERS_2_39_port, 
      REGISTERS_2_38_port, REGISTERS_2_37_port, REGISTERS_2_36_port, 
      REGISTERS_2_35_port, REGISTERS_2_34_port, REGISTERS_2_33_port, 
      REGISTERS_2_32_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_63_port, REGISTERS_3_62_port, REGISTERS_3_61_port, 
      REGISTERS_3_60_port, REGISTERS_3_59_port, REGISTERS_3_58_port, 
      REGISTERS_3_57_port, REGISTERS_3_56_port, REGISTERS_3_55_port, 
      REGISTERS_3_54_port, REGISTERS_3_53_port, REGISTERS_3_52_port, 
      REGISTERS_3_51_port, REGISTERS_3_50_port, REGISTERS_3_49_port, 
      REGISTERS_3_48_port, REGISTERS_3_47_port, REGISTERS_3_46_port, 
      REGISTERS_3_45_port, REGISTERS_3_44_port, REGISTERS_3_43_port, 
      REGISTERS_3_42_port, REGISTERS_3_41_port, REGISTERS_3_40_port, 
      REGISTERS_3_39_port, REGISTERS_3_38_port, REGISTERS_3_37_port, 
      REGISTERS_3_36_port, REGISTERS_3_35_port, REGISTERS_3_34_port, 
      REGISTERS_3_33_port, REGISTERS_3_32_port, REGISTERS_3_31_port, 
      REGISTERS_3_30_port, REGISTERS_3_29_port, REGISTERS_3_28_port, 
      REGISTERS_3_27_port, REGISTERS_3_26_port, REGISTERS_3_25_port, 
      REGISTERS_3_24_port, REGISTERS_3_23_port, REGISTERS_3_22_port, 
      REGISTERS_3_21_port, REGISTERS_3_20_port, REGISTERS_3_19_port, 
      REGISTERS_3_18_port, REGISTERS_3_17_port, REGISTERS_3_16_port, 
      REGISTERS_3_15_port, REGISTERS_3_14_port, REGISTERS_3_13_port, 
      REGISTERS_3_12_port, REGISTERS_3_11_port, REGISTERS_3_10_port, 
      REGISTERS_3_9_port, REGISTERS_3_8_port, REGISTERS_3_7_port, 
      REGISTERS_3_6_port, REGISTERS_3_5_port, REGISTERS_3_4_port, 
      REGISTERS_3_3_port, REGISTERS_3_2_port, REGISTERS_3_1_port, 
      REGISTERS_3_0_port, REGISTERS_4_63_port, REGISTERS_4_62_port, 
      REGISTERS_4_61_port, REGISTERS_4_60_port, REGISTERS_4_59_port, 
      REGISTERS_4_58_port, REGISTERS_4_57_port, REGISTERS_4_56_port, 
      REGISTERS_4_55_port, REGISTERS_4_54_port, REGISTERS_4_53_port, 
      REGISTERS_4_52_port, REGISTERS_4_51_port, REGISTERS_4_50_port, 
      REGISTERS_4_49_port, REGISTERS_4_48_port, REGISTERS_4_47_port, 
      REGISTERS_4_46_port, REGISTERS_4_45_port, REGISTERS_4_44_port, 
      REGISTERS_4_43_port, REGISTERS_4_42_port, REGISTERS_4_41_port, 
      REGISTERS_4_40_port, REGISTERS_4_39_port, REGISTERS_4_38_port, 
      REGISTERS_4_37_port, REGISTERS_4_36_port, REGISTERS_4_35_port, 
      REGISTERS_4_34_port, REGISTERS_4_33_port, REGISTERS_4_32_port, 
      REGISTERS_4_31_port, REGISTERS_4_30_port, REGISTERS_4_29_port, 
      REGISTERS_4_28_port, REGISTERS_4_27_port, REGISTERS_4_26_port, 
      REGISTERS_4_25_port, REGISTERS_4_24_port, REGISTERS_4_23_port, 
      REGISTERS_4_22_port, REGISTERS_4_21_port, REGISTERS_4_20_port, 
      REGISTERS_4_19_port, REGISTERS_4_18_port, REGISTERS_4_17_port, 
      REGISTERS_4_16_port, REGISTERS_4_15_port, REGISTERS_4_14_port, 
      REGISTERS_4_13_port, REGISTERS_4_12_port, REGISTERS_4_11_port, 
      REGISTERS_4_10_port, REGISTERS_4_9_port, REGISTERS_4_8_port, 
      REGISTERS_4_7_port, REGISTERS_4_6_port, REGISTERS_4_5_port, 
      REGISTERS_4_4_port, REGISTERS_4_3_port, REGISTERS_4_2_port, 
      REGISTERS_4_1_port, REGISTERS_4_0_port, REGISTERS_5_63_port, 
      REGISTERS_5_62_port, REGISTERS_5_61_port, REGISTERS_5_60_port, 
      REGISTERS_5_59_port, REGISTERS_5_58_port, REGISTERS_5_57_port, 
      REGISTERS_5_56_port, REGISTERS_5_55_port, REGISTERS_5_54_port, 
      REGISTERS_5_53_port, REGISTERS_5_52_port, REGISTERS_5_51_port, 
      REGISTERS_5_50_port, REGISTERS_5_49_port, REGISTERS_5_48_port, 
      REGISTERS_5_47_port, REGISTERS_5_46_port, REGISTERS_5_45_port, 
      REGISTERS_5_44_port, REGISTERS_5_43_port, REGISTERS_5_42_port, 
      REGISTERS_5_41_port, REGISTERS_5_40_port, REGISTERS_5_39_port, 
      REGISTERS_5_38_port, REGISTERS_5_37_port, REGISTERS_5_36_port, 
      REGISTERS_5_35_port, REGISTERS_5_34_port, REGISTERS_5_33_port, 
      REGISTERS_5_32_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_63_port, REGISTERS_6_62_port, REGISTERS_6_61_port, 
      REGISTERS_6_60_port, REGISTERS_6_59_port, REGISTERS_6_58_port, 
      REGISTERS_6_57_port, REGISTERS_6_56_port, REGISTERS_6_55_port, 
      REGISTERS_6_54_port, REGISTERS_6_53_port, REGISTERS_6_52_port, 
      REGISTERS_6_51_port, REGISTERS_6_50_port, REGISTERS_6_49_port, 
      REGISTERS_6_48_port, REGISTERS_6_47_port, REGISTERS_6_46_port, 
      REGISTERS_6_45_port, REGISTERS_6_44_port, REGISTERS_6_43_port, 
      REGISTERS_6_42_port, REGISTERS_6_41_port, REGISTERS_6_40_port, 
      REGISTERS_6_39_port, REGISTERS_6_38_port, REGISTERS_6_37_port, 
      REGISTERS_6_36_port, REGISTERS_6_35_port, REGISTERS_6_34_port, 
      REGISTERS_6_33_port, REGISTERS_6_32_port, REGISTERS_6_31_port, 
      REGISTERS_6_30_port, REGISTERS_6_29_port, REGISTERS_6_28_port, 
      REGISTERS_6_27_port, REGISTERS_6_26_port, REGISTERS_6_25_port, 
      REGISTERS_6_24_port, REGISTERS_6_23_port, REGISTERS_6_22_port, 
      REGISTERS_6_21_port, REGISTERS_6_20_port, REGISTERS_6_19_port, 
      REGISTERS_6_18_port, REGISTERS_6_17_port, REGISTERS_6_16_port, 
      REGISTERS_6_15_port, REGISTERS_6_14_port, REGISTERS_6_13_port, 
      REGISTERS_6_12_port, REGISTERS_6_11_port, REGISTERS_6_10_port, 
      REGISTERS_6_9_port, REGISTERS_6_8_port, REGISTERS_6_7_port, 
      REGISTERS_6_6_port, REGISTERS_6_5_port, REGISTERS_6_4_port, 
      REGISTERS_6_3_port, REGISTERS_6_2_port, REGISTERS_6_1_port, 
      REGISTERS_6_0_port, REGISTERS_7_63_port, REGISTERS_7_62_port, 
      REGISTERS_7_61_port, REGISTERS_7_60_port, REGISTERS_7_59_port, 
      REGISTERS_7_58_port, REGISTERS_7_57_port, REGISTERS_7_56_port, 
      REGISTERS_7_55_port, REGISTERS_7_54_port, REGISTERS_7_53_port, 
      REGISTERS_7_52_port, REGISTERS_7_51_port, REGISTERS_7_50_port, 
      REGISTERS_7_49_port, REGISTERS_7_48_port, REGISTERS_7_47_port, 
      REGISTERS_7_46_port, REGISTERS_7_45_port, REGISTERS_7_44_port, 
      REGISTERS_7_43_port, REGISTERS_7_42_port, REGISTERS_7_41_port, 
      REGISTERS_7_40_port, REGISTERS_7_39_port, REGISTERS_7_38_port, 
      REGISTERS_7_37_port, REGISTERS_7_36_port, REGISTERS_7_35_port, 
      REGISTERS_7_34_port, REGISTERS_7_33_port, REGISTERS_7_32_port, 
      REGISTERS_7_31_port, REGISTERS_7_30_port, REGISTERS_7_29_port, 
      REGISTERS_7_28_port, REGISTERS_7_27_port, REGISTERS_7_26_port, 
      REGISTERS_7_25_port, REGISTERS_7_24_port, REGISTERS_7_23_port, 
      REGISTERS_7_22_port, REGISTERS_7_21_port, REGISTERS_7_20_port, 
      REGISTERS_7_19_port, REGISTERS_7_18_port, REGISTERS_7_17_port, 
      REGISTERS_7_16_port, REGISTERS_7_15_port, REGISTERS_7_14_port, 
      REGISTERS_7_13_port, REGISTERS_7_12_port, REGISTERS_7_11_port, 
      REGISTERS_7_10_port, REGISTERS_7_9_port, REGISTERS_7_8_port, 
      REGISTERS_7_7_port, REGISTERS_7_6_port, REGISTERS_7_5_port, 
      REGISTERS_7_4_port, REGISTERS_7_3_port, REGISTERS_7_2_port, 
      REGISTERS_7_1_port, REGISTERS_7_0_port, REGISTERS_8_63_port, 
      REGISTERS_8_62_port, REGISTERS_8_61_port, REGISTERS_8_60_port, 
      REGISTERS_8_59_port, REGISTERS_8_58_port, REGISTERS_8_57_port, 
      REGISTERS_8_56_port, REGISTERS_8_55_port, REGISTERS_8_54_port, 
      REGISTERS_8_53_port, REGISTERS_8_52_port, REGISTERS_8_51_port, 
      REGISTERS_8_50_port, REGISTERS_8_49_port, REGISTERS_8_48_port, 
      REGISTERS_8_47_port, REGISTERS_8_46_port, REGISTERS_8_45_port, 
      REGISTERS_8_44_port, REGISTERS_8_43_port, REGISTERS_8_42_port, 
      REGISTERS_8_41_port, REGISTERS_8_40_port, REGISTERS_8_39_port, 
      REGISTERS_8_38_port, REGISTERS_8_37_port, REGISTERS_8_36_port, 
      REGISTERS_8_35_port, REGISTERS_8_34_port, REGISTERS_8_33_port, 
      REGISTERS_8_32_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_63_port, REGISTERS_9_62_port, REGISTERS_9_61_port, 
      REGISTERS_9_60_port, REGISTERS_9_59_port, REGISTERS_9_58_port, 
      REGISTERS_9_57_port, REGISTERS_9_56_port, REGISTERS_9_55_port, 
      REGISTERS_9_54_port, REGISTERS_9_53_port, REGISTERS_9_52_port, 
      REGISTERS_9_51_port, REGISTERS_9_50_port, REGISTERS_9_49_port, 
      REGISTERS_9_48_port, REGISTERS_9_47_port, REGISTERS_9_46_port, 
      REGISTERS_9_45_port, REGISTERS_9_44_port, REGISTERS_9_43_port, 
      REGISTERS_9_42_port, REGISTERS_9_41_port, REGISTERS_9_40_port, 
      REGISTERS_9_39_port, REGISTERS_9_38_port, REGISTERS_9_37_port, 
      REGISTERS_9_36_port, REGISTERS_9_35_port, REGISTERS_9_34_port, 
      REGISTERS_9_33_port, REGISTERS_9_32_port, REGISTERS_9_31_port, 
      REGISTERS_9_30_port, REGISTERS_9_29_port, REGISTERS_9_28_port, 
      REGISTERS_9_27_port, REGISTERS_9_26_port, REGISTERS_9_25_port, 
      REGISTERS_9_24_port, REGISTERS_9_23_port, REGISTERS_9_22_port, 
      REGISTERS_9_21_port, REGISTERS_9_20_port, REGISTERS_9_19_port, 
      REGISTERS_9_18_port, REGISTERS_9_17_port, REGISTERS_9_16_port, 
      REGISTERS_9_15_port, REGISTERS_9_14_port, REGISTERS_9_13_port, 
      REGISTERS_9_12_port, REGISTERS_9_11_port, REGISTERS_9_10_port, 
      REGISTERS_9_9_port, REGISTERS_9_8_port, REGISTERS_9_7_port, 
      REGISTERS_9_6_port, REGISTERS_9_5_port, REGISTERS_9_4_port, 
      REGISTERS_9_3_port, REGISTERS_9_2_port, REGISTERS_9_1_port, 
      REGISTERS_9_0_port, REGISTERS_10_63_port, REGISTERS_10_62_port, 
      REGISTERS_10_61_port, REGISTERS_10_60_port, REGISTERS_10_59_port, 
      REGISTERS_10_58_port, REGISTERS_10_57_port, REGISTERS_10_56_port, 
      REGISTERS_10_55_port, REGISTERS_10_54_port, REGISTERS_10_53_port, 
      REGISTERS_10_52_port, REGISTERS_10_51_port, REGISTERS_10_50_port, 
      REGISTERS_10_49_port, REGISTERS_10_48_port, REGISTERS_10_47_port, 
      REGISTERS_10_46_port, REGISTERS_10_45_port, REGISTERS_10_44_port, 
      REGISTERS_10_43_port, REGISTERS_10_42_port, REGISTERS_10_41_port, 
      REGISTERS_10_40_port, REGISTERS_10_39_port, REGISTERS_10_38_port, 
      REGISTERS_10_37_port, REGISTERS_10_36_port, REGISTERS_10_35_port, 
      REGISTERS_10_34_port, REGISTERS_10_33_port, REGISTERS_10_32_port, 
      REGISTERS_10_31_port, REGISTERS_10_30_port, REGISTERS_10_29_port, 
      REGISTERS_10_28_port, REGISTERS_10_27_port, REGISTERS_10_26_port, 
      REGISTERS_10_25_port, REGISTERS_10_24_port, REGISTERS_10_23_port, 
      REGISTERS_10_22_port, REGISTERS_10_21_port, REGISTERS_10_20_port, 
      REGISTERS_10_19_port, REGISTERS_10_18_port, REGISTERS_10_17_port, 
      REGISTERS_10_16_port, REGISTERS_10_15_port, REGISTERS_10_14_port, 
      REGISTERS_10_13_port, REGISTERS_10_12_port, REGISTERS_10_11_port, 
      REGISTERS_10_10_port, REGISTERS_10_9_port, REGISTERS_10_8_port, 
      REGISTERS_10_7_port, REGISTERS_10_6_port, REGISTERS_10_5_port, 
      REGISTERS_10_4_port, REGISTERS_10_3_port, REGISTERS_10_2_port, 
      REGISTERS_10_1_port, REGISTERS_10_0_port, REGISTERS_11_63_port, 
      REGISTERS_11_62_port, REGISTERS_11_61_port, REGISTERS_11_60_port, 
      REGISTERS_11_59_port, REGISTERS_11_58_port, REGISTERS_11_57_port, 
      REGISTERS_11_56_port, REGISTERS_11_55_port, REGISTERS_11_54_port, 
      REGISTERS_11_53_port, REGISTERS_11_52_port, REGISTERS_11_51_port, 
      REGISTERS_11_50_port, REGISTERS_11_49_port, REGISTERS_11_48_port, 
      REGISTERS_11_47_port, REGISTERS_11_46_port, REGISTERS_11_45_port, 
      REGISTERS_11_44_port, REGISTERS_11_43_port, REGISTERS_11_42_port, 
      REGISTERS_11_41_port, REGISTERS_11_40_port, REGISTERS_11_39_port, 
      REGISTERS_11_38_port, REGISTERS_11_37_port, REGISTERS_11_36_port, 
      REGISTERS_11_35_port, REGISTERS_11_34_port, REGISTERS_11_33_port, 
      REGISTERS_11_32_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_63_port, REGISTERS_12_62_port, REGISTERS_12_61_port, 
      REGISTERS_12_60_port, REGISTERS_12_59_port, REGISTERS_12_58_port, 
      REGISTERS_12_57_port, REGISTERS_12_56_port, REGISTERS_12_55_port, 
      REGISTERS_12_54_port, REGISTERS_12_53_port, REGISTERS_12_52_port, 
      REGISTERS_12_51_port, REGISTERS_12_50_port, REGISTERS_12_49_port, 
      REGISTERS_12_48_port, REGISTERS_12_47_port, REGISTERS_12_46_port, 
      REGISTERS_12_45_port, REGISTERS_12_44_port, REGISTERS_12_43_port, 
      REGISTERS_12_42_port, REGISTERS_12_41_port, REGISTERS_12_40_port, 
      REGISTERS_12_39_port, REGISTERS_12_38_port, REGISTERS_12_37_port, 
      REGISTERS_12_36_port, REGISTERS_12_35_port, REGISTERS_12_34_port, 
      REGISTERS_12_33_port, REGISTERS_12_32_port, REGISTERS_12_31_port, 
      REGISTERS_12_30_port, REGISTERS_12_29_port, REGISTERS_12_28_port, 
      REGISTERS_12_27_port, REGISTERS_12_26_port, REGISTERS_12_25_port, 
      REGISTERS_12_24_port, REGISTERS_12_23_port, REGISTERS_12_22_port, 
      REGISTERS_12_21_port, REGISTERS_12_20_port, REGISTERS_12_19_port, 
      REGISTERS_12_18_port, REGISTERS_12_17_port, REGISTERS_12_16_port, 
      REGISTERS_12_15_port, REGISTERS_12_14_port, REGISTERS_12_13_port, 
      REGISTERS_12_12_port, REGISTERS_12_11_port, REGISTERS_12_10_port, 
      REGISTERS_12_9_port, REGISTERS_12_8_port, REGISTERS_12_7_port, 
      REGISTERS_12_6_port, REGISTERS_12_5_port, REGISTERS_12_4_port, 
      REGISTERS_12_3_port, REGISTERS_12_2_port, REGISTERS_12_1_port, 
      REGISTERS_12_0_port, REGISTERS_13_63_port, REGISTERS_13_62_port, 
      REGISTERS_13_61_port, REGISTERS_13_60_port, REGISTERS_13_59_port, 
      REGISTERS_13_58_port, REGISTERS_13_57_port, REGISTERS_13_56_port, 
      REGISTERS_13_55_port, REGISTERS_13_54_port, REGISTERS_13_53_port, 
      REGISTERS_13_52_port, REGISTERS_13_51_port, REGISTERS_13_50_port, 
      REGISTERS_13_49_port, REGISTERS_13_48_port, REGISTERS_13_47_port, 
      REGISTERS_13_46_port, REGISTERS_13_45_port, REGISTERS_13_44_port, 
      REGISTERS_13_43_port, REGISTERS_13_42_port, REGISTERS_13_41_port, 
      REGISTERS_13_40_port, REGISTERS_13_39_port, REGISTERS_13_38_port, 
      REGISTERS_13_37_port, REGISTERS_13_36_port, REGISTERS_13_35_port, 
      REGISTERS_13_34_port, REGISTERS_13_33_port, REGISTERS_13_32_port, 
      REGISTERS_13_31_port, REGISTERS_13_30_port, REGISTERS_13_29_port, 
      REGISTERS_13_28_port, REGISTERS_13_27_port, REGISTERS_13_26_port, 
      REGISTERS_13_25_port, REGISTERS_13_24_port, REGISTERS_13_23_port, 
      REGISTERS_13_22_port, REGISTERS_13_21_port, REGISTERS_13_20_port, 
      REGISTERS_13_19_port, REGISTERS_13_18_port, REGISTERS_13_17_port, 
      REGISTERS_13_16_port, REGISTERS_13_15_port, REGISTERS_13_14_port, 
      REGISTERS_13_13_port, REGISTERS_13_12_port, REGISTERS_13_11_port, 
      REGISTERS_13_10_port, REGISTERS_13_9_port, REGISTERS_13_8_port, 
      REGISTERS_13_7_port, REGISTERS_13_6_port, REGISTERS_13_5_port, 
      REGISTERS_13_4_port, REGISTERS_13_3_port, REGISTERS_13_2_port, 
      REGISTERS_13_1_port, REGISTERS_13_0_port, REGISTERS_14_63_port, 
      REGISTERS_14_62_port, REGISTERS_14_61_port, REGISTERS_14_60_port, 
      REGISTERS_14_59_port, REGISTERS_14_58_port, REGISTERS_14_57_port, 
      REGISTERS_14_56_port, REGISTERS_14_55_port, REGISTERS_14_54_port, 
      REGISTERS_14_53_port, REGISTERS_14_52_port, REGISTERS_14_51_port, 
      REGISTERS_14_50_port, REGISTERS_14_49_port, REGISTERS_14_48_port, 
      REGISTERS_14_47_port, REGISTERS_14_46_port, REGISTERS_14_45_port, 
      REGISTERS_14_44_port, REGISTERS_14_43_port, REGISTERS_14_42_port, 
      REGISTERS_14_41_port, REGISTERS_14_40_port, REGISTERS_14_39_port, 
      REGISTERS_14_38_port, REGISTERS_14_37_port, REGISTERS_14_36_port, 
      REGISTERS_14_35_port, REGISTERS_14_34_port, REGISTERS_14_33_port, 
      REGISTERS_14_32_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_63_port, REGISTERS_15_62_port, REGISTERS_15_61_port, 
      REGISTERS_15_60_port, REGISTERS_15_59_port, REGISTERS_15_58_port, 
      REGISTERS_15_57_port, REGISTERS_15_56_port, REGISTERS_15_55_port, 
      REGISTERS_15_54_port, REGISTERS_15_53_port, REGISTERS_15_52_port, 
      REGISTERS_15_51_port, REGISTERS_15_50_port, REGISTERS_15_49_port, 
      REGISTERS_15_48_port, REGISTERS_15_47_port, REGISTERS_15_46_port, 
      REGISTERS_15_45_port, REGISTERS_15_44_port, REGISTERS_15_43_port, 
      REGISTERS_15_42_port, REGISTERS_15_41_port, REGISTERS_15_40_port, 
      REGISTERS_15_39_port, REGISTERS_15_38_port, REGISTERS_15_37_port, 
      REGISTERS_15_36_port, REGISTERS_15_35_port, REGISTERS_15_34_port, 
      REGISTERS_15_33_port, REGISTERS_15_32_port, REGISTERS_15_31_port, 
      REGISTERS_15_30_port, REGISTERS_15_29_port, REGISTERS_15_28_port, 
      REGISTERS_15_27_port, REGISTERS_15_26_port, REGISTERS_15_25_port, 
      REGISTERS_15_24_port, REGISTERS_15_23_port, REGISTERS_15_22_port, 
      REGISTERS_15_21_port, REGISTERS_15_20_port, REGISTERS_15_19_port, 
      REGISTERS_15_18_port, REGISTERS_15_17_port, REGISTERS_15_16_port, 
      REGISTERS_15_15_port, REGISTERS_15_14_port, REGISTERS_15_13_port, 
      REGISTERS_15_12_port, REGISTERS_15_11_port, REGISTERS_15_10_port, 
      REGISTERS_15_9_port, REGISTERS_15_8_port, REGISTERS_15_7_port, 
      REGISTERS_15_6_port, REGISTERS_15_5_port, REGISTERS_15_4_port, 
      REGISTERS_15_3_port, REGISTERS_15_2_port, REGISTERS_15_1_port, 
      REGISTERS_15_0_port, REGISTERS_16_63_port, REGISTERS_16_62_port, 
      REGISTERS_16_61_port, REGISTERS_16_60_port, REGISTERS_16_59_port, 
      REGISTERS_16_58_port, REGISTERS_16_57_port, REGISTERS_16_56_port, 
      REGISTERS_16_55_port, REGISTERS_16_54_port, REGISTERS_16_53_port, 
      REGISTERS_16_52_port, REGISTERS_16_51_port, REGISTERS_16_50_port, 
      REGISTERS_16_49_port, REGISTERS_16_48_port, REGISTERS_16_47_port, 
      REGISTERS_16_46_port, REGISTERS_16_45_port, REGISTERS_16_44_port, 
      REGISTERS_16_43_port, REGISTERS_16_42_port, REGISTERS_16_41_port, 
      REGISTERS_16_40_port, REGISTERS_16_39_port, REGISTERS_16_38_port, 
      REGISTERS_16_37_port, REGISTERS_16_36_port, REGISTERS_16_35_port, 
      REGISTERS_16_34_port, REGISTERS_16_33_port, REGISTERS_16_32_port, 
      REGISTERS_16_31_port, REGISTERS_16_30_port, REGISTERS_16_29_port, 
      REGISTERS_16_28_port, REGISTERS_16_27_port, REGISTERS_16_26_port, 
      REGISTERS_16_25_port, REGISTERS_16_24_port, REGISTERS_16_23_port, 
      REGISTERS_16_22_port, REGISTERS_16_21_port, REGISTERS_16_20_port, 
      REGISTERS_16_19_port, REGISTERS_16_18_port, REGISTERS_16_17_port, 
      REGISTERS_16_16_port, REGISTERS_16_15_port, REGISTERS_16_14_port, 
      REGISTERS_16_13_port, REGISTERS_16_12_port, REGISTERS_16_11_port, 
      REGISTERS_16_10_port, REGISTERS_16_9_port, REGISTERS_16_8_port, 
      REGISTERS_16_7_port, REGISTERS_16_6_port, REGISTERS_16_5_port, 
      REGISTERS_16_4_port, REGISTERS_16_3_port, REGISTERS_16_2_port, 
      REGISTERS_16_1_port, REGISTERS_16_0_port, REGISTERS_17_63_port, 
      REGISTERS_17_62_port, REGISTERS_17_61_port, REGISTERS_17_60_port, 
      REGISTERS_17_59_port, REGISTERS_17_58_port, REGISTERS_17_57_port, 
      REGISTERS_17_56_port, REGISTERS_17_55_port, REGISTERS_17_54_port, 
      REGISTERS_17_53_port, REGISTERS_17_52_port, REGISTERS_17_51_port, 
      REGISTERS_17_50_port, REGISTERS_17_49_port, REGISTERS_17_48_port, 
      REGISTERS_17_47_port, REGISTERS_17_46_port, REGISTERS_17_45_port, 
      REGISTERS_17_44_port, REGISTERS_17_43_port, REGISTERS_17_42_port, 
      REGISTERS_17_41_port, REGISTERS_17_40_port, REGISTERS_17_39_port, 
      REGISTERS_17_38_port, REGISTERS_17_37_port, REGISTERS_17_36_port, 
      REGISTERS_17_35_port, REGISTERS_17_34_port, REGISTERS_17_33_port, 
      REGISTERS_17_32_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_63_port, REGISTERS_18_62_port, REGISTERS_18_61_port, 
      REGISTERS_18_60_port, REGISTERS_18_59_port, REGISTERS_18_58_port, 
      REGISTERS_18_57_port, REGISTERS_18_56_port, REGISTERS_18_55_port, 
      REGISTERS_18_54_port, REGISTERS_18_53_port, REGISTERS_18_52_port, 
      REGISTERS_18_51_port, REGISTERS_18_50_port, REGISTERS_18_49_port, 
      REGISTERS_18_48_port, REGISTERS_18_47_port, REGISTERS_18_46_port, 
      REGISTERS_18_45_port, REGISTERS_18_44_port, REGISTERS_18_43_port, 
      REGISTERS_18_42_port, REGISTERS_18_41_port, REGISTERS_18_40_port, 
      REGISTERS_18_39_port, REGISTERS_18_38_port, REGISTERS_18_37_port, 
      REGISTERS_18_36_port, REGISTERS_18_35_port, REGISTERS_18_34_port, 
      REGISTERS_18_33_port, REGISTERS_18_32_port, REGISTERS_18_31_port, 
      REGISTERS_18_30_port, REGISTERS_18_29_port, REGISTERS_18_28_port, 
      REGISTERS_18_27_port, REGISTERS_18_26_port, REGISTERS_18_25_port, 
      REGISTERS_18_24_port, REGISTERS_18_23_port, REGISTERS_18_22_port, 
      REGISTERS_18_21_port, REGISTERS_18_20_port, REGISTERS_18_19_port, 
      REGISTERS_18_18_port, REGISTERS_18_17_port, REGISTERS_18_16_port, 
      REGISTERS_18_15_port, REGISTERS_18_14_port, REGISTERS_18_13_port, 
      REGISTERS_18_12_port, REGISTERS_18_11_port, REGISTERS_18_10_port, 
      REGISTERS_18_9_port, REGISTERS_18_8_port, REGISTERS_18_7_port, 
      REGISTERS_18_6_port, REGISTERS_18_5_port, REGISTERS_18_4_port, 
      REGISTERS_18_3_port, REGISTERS_18_2_port, REGISTERS_18_1_port, 
      REGISTERS_18_0_port, REGISTERS_19_63_port, REGISTERS_19_62_port, 
      REGISTERS_19_61_port, REGISTERS_19_60_port, REGISTERS_19_59_port, 
      REGISTERS_19_58_port, REGISTERS_19_57_port, REGISTERS_19_56_port, 
      REGISTERS_19_55_port, REGISTERS_19_54_port, REGISTERS_19_53_port, 
      REGISTERS_19_52_port, REGISTERS_19_51_port, REGISTERS_19_50_port, 
      REGISTERS_19_49_port, REGISTERS_19_48_port, REGISTERS_19_47_port, 
      REGISTERS_19_46_port, REGISTERS_19_45_port, REGISTERS_19_44_port, 
      REGISTERS_19_43_port, REGISTERS_19_42_port, REGISTERS_19_41_port, 
      REGISTERS_19_40_port, REGISTERS_19_39_port, REGISTERS_19_38_port, 
      REGISTERS_19_37_port, REGISTERS_19_36_port, REGISTERS_19_35_port, 
      REGISTERS_19_34_port, REGISTERS_19_33_port, REGISTERS_19_32_port, 
      REGISTERS_19_31_port, REGISTERS_19_30_port, REGISTERS_19_29_port, 
      REGISTERS_19_28_port, REGISTERS_19_27_port, REGISTERS_19_26_port, 
      REGISTERS_19_25_port, REGISTERS_19_24_port, REGISTERS_19_23_port, 
      REGISTERS_19_22_port, REGISTERS_19_21_port, REGISTERS_19_20_port, 
      REGISTERS_19_19_port, REGISTERS_19_18_port, REGISTERS_19_17_port, 
      REGISTERS_19_16_port, REGISTERS_19_15_port, REGISTERS_19_14_port, 
      REGISTERS_19_13_port, REGISTERS_19_12_port, REGISTERS_19_11_port, 
      REGISTERS_19_10_port, REGISTERS_19_9_port, REGISTERS_19_8_port, 
      REGISTERS_19_7_port, REGISTERS_19_6_port, REGISTERS_19_5_port, 
      REGISTERS_19_4_port, REGISTERS_19_3_port, REGISTERS_19_2_port, 
      REGISTERS_19_1_port, REGISTERS_19_0_port, REGISTERS_20_63_port, 
      REGISTERS_20_62_port, REGISTERS_20_61_port, REGISTERS_20_60_port, 
      REGISTERS_20_59_port, REGISTERS_20_58_port, REGISTERS_20_57_port, 
      REGISTERS_20_56_port, REGISTERS_20_55_port, REGISTERS_20_54_port, 
      REGISTERS_20_53_port, REGISTERS_20_52_port, REGISTERS_20_51_port, 
      REGISTERS_20_50_port, REGISTERS_20_49_port, REGISTERS_20_48_port, 
      REGISTERS_20_47_port, REGISTERS_20_46_port, REGISTERS_20_45_port, 
      REGISTERS_20_44_port, REGISTERS_20_43_port, REGISTERS_20_42_port, 
      REGISTERS_20_41_port, REGISTERS_20_40_port, REGISTERS_20_39_port, 
      REGISTERS_20_38_port, REGISTERS_20_37_port, REGISTERS_20_36_port, 
      REGISTERS_20_35_port, REGISTERS_20_34_port, REGISTERS_20_33_port, 
      REGISTERS_20_32_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_63_port, REGISTERS_21_62_port, REGISTERS_21_61_port, 
      REGISTERS_21_60_port, REGISTERS_21_59_port, REGISTERS_21_58_port, 
      REGISTERS_21_57_port, REGISTERS_21_56_port, REGISTERS_21_55_port, 
      REGISTERS_21_54_port, REGISTERS_21_53_port, REGISTERS_21_52_port, 
      REGISTERS_21_51_port, REGISTERS_21_50_port, REGISTERS_21_49_port, 
      REGISTERS_21_48_port, REGISTERS_21_47_port, REGISTERS_21_46_port, 
      REGISTERS_21_45_port, REGISTERS_21_44_port, REGISTERS_21_43_port, 
      REGISTERS_21_42_port, REGISTERS_21_41_port, REGISTERS_21_40_port, 
      REGISTERS_21_39_port, REGISTERS_21_38_port, REGISTERS_21_37_port, 
      REGISTERS_21_36_port, REGISTERS_21_35_port, REGISTERS_21_34_port, 
      REGISTERS_21_33_port, REGISTERS_21_32_port, REGISTERS_21_31_port, 
      REGISTERS_21_30_port, REGISTERS_21_29_port, REGISTERS_21_28_port, 
      REGISTERS_21_27_port, REGISTERS_21_26_port, REGISTERS_21_25_port, 
      REGISTERS_21_24_port, REGISTERS_21_23_port, REGISTERS_21_22_port, 
      REGISTERS_21_21_port, REGISTERS_21_20_port, REGISTERS_21_19_port, 
      REGISTERS_21_18_port, REGISTERS_21_17_port, REGISTERS_21_16_port, 
      REGISTERS_21_15_port, REGISTERS_21_14_port, REGISTERS_21_13_port, 
      REGISTERS_21_12_port, REGISTERS_21_11_port, REGISTERS_21_10_port, 
      REGISTERS_21_9_port, REGISTERS_21_8_port, REGISTERS_21_7_port, 
      REGISTERS_21_6_port, REGISTERS_21_5_port, REGISTERS_21_4_port, 
      REGISTERS_21_3_port, REGISTERS_21_2_port, REGISTERS_21_1_port, 
      REGISTERS_21_0_port, REGISTERS_22_63_port, REGISTERS_22_62_port, 
      REGISTERS_22_61_port, REGISTERS_22_60_port, REGISTERS_22_59_port, 
      REGISTERS_22_58_port, REGISTERS_22_57_port, REGISTERS_22_56_port, 
      REGISTERS_22_55_port, REGISTERS_22_54_port, REGISTERS_22_53_port, 
      REGISTERS_22_52_port, REGISTERS_22_51_port, REGISTERS_22_50_port, 
      REGISTERS_22_49_port, REGISTERS_22_48_port, REGISTERS_22_47_port, 
      REGISTERS_22_46_port, REGISTERS_22_45_port, REGISTERS_22_44_port, 
      REGISTERS_22_43_port, REGISTERS_22_42_port, REGISTERS_22_41_port, 
      REGISTERS_22_40_port, REGISTERS_22_39_port, REGISTERS_22_38_port, 
      REGISTERS_22_37_port, REGISTERS_22_36_port, REGISTERS_22_35_port, 
      REGISTERS_22_34_port, REGISTERS_22_33_port, REGISTERS_22_32_port, 
      REGISTERS_22_31_port, REGISTERS_22_30_port, REGISTERS_22_29_port, 
      REGISTERS_22_28_port, REGISTERS_22_27_port, REGISTERS_22_26_port, 
      REGISTERS_22_25_port, REGISTERS_22_24_port, REGISTERS_22_23_port, 
      REGISTERS_22_22_port, REGISTERS_22_21_port, REGISTERS_22_20_port, 
      REGISTERS_22_19_port, REGISTERS_22_18_port, REGISTERS_22_17_port, 
      REGISTERS_22_16_port, REGISTERS_22_15_port, REGISTERS_22_14_port, 
      REGISTERS_22_13_port, REGISTERS_22_12_port, REGISTERS_22_11_port, 
      REGISTERS_22_10_port, REGISTERS_22_9_port, REGISTERS_22_8_port, 
      REGISTERS_22_7_port, REGISTERS_22_6_port, REGISTERS_22_5_port, 
      REGISTERS_22_4_port, REGISTERS_22_3_port, REGISTERS_22_2_port, 
      REGISTERS_22_1_port, REGISTERS_22_0_port, REGISTERS_23_63_port, 
      REGISTERS_23_62_port, REGISTERS_23_61_port, REGISTERS_23_60_port, 
      REGISTERS_23_59_port, REGISTERS_23_58_port, REGISTERS_23_57_port, 
      REGISTERS_23_56_port, REGISTERS_23_55_port, REGISTERS_23_54_port, 
      REGISTERS_23_53_port, REGISTERS_23_52_port, REGISTERS_23_51_port, 
      REGISTERS_23_50_port, REGISTERS_23_49_port, REGISTERS_23_48_port, 
      REGISTERS_23_47_port, REGISTERS_23_46_port, REGISTERS_23_45_port, 
      REGISTERS_23_44_port, REGISTERS_23_43_port, REGISTERS_23_42_port, 
      REGISTERS_23_41_port, REGISTERS_23_40_port, REGISTERS_23_39_port, 
      REGISTERS_23_38_port, REGISTERS_23_37_port, REGISTERS_23_36_port, 
      REGISTERS_23_35_port, REGISTERS_23_34_port, REGISTERS_23_33_port, 
      REGISTERS_23_32_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_63_port, REGISTERS_24_62_port, REGISTERS_24_61_port, 
      REGISTERS_24_60_port, REGISTERS_24_59_port, REGISTERS_24_58_port, 
      REGISTERS_24_57_port, REGISTERS_24_56_port, REGISTERS_24_55_port, 
      REGISTERS_24_54_port, REGISTERS_24_53_port, REGISTERS_24_52_port, 
      REGISTERS_24_51_port, REGISTERS_24_50_port, REGISTERS_24_49_port, 
      REGISTERS_24_48_port, REGISTERS_24_47_port, REGISTERS_24_46_port, 
      REGISTERS_24_45_port, REGISTERS_24_44_port, REGISTERS_24_43_port, 
      REGISTERS_24_42_port, REGISTERS_24_41_port, REGISTERS_24_40_port, 
      REGISTERS_24_39_port, REGISTERS_24_38_port, REGISTERS_24_37_port, 
      REGISTERS_24_36_port, REGISTERS_24_35_port, REGISTERS_24_34_port, 
      REGISTERS_24_33_port, REGISTERS_24_32_port, REGISTERS_24_31_port, 
      REGISTERS_24_30_port, REGISTERS_24_29_port, REGISTERS_24_28_port, 
      REGISTERS_24_27_port, REGISTERS_24_26_port, REGISTERS_24_25_port, 
      REGISTERS_24_24_port, REGISTERS_24_23_port, REGISTERS_24_22_port, 
      REGISTERS_24_21_port, REGISTERS_24_20_port, REGISTERS_24_19_port, 
      REGISTERS_24_18_port, REGISTERS_24_17_port, REGISTERS_24_16_port, 
      REGISTERS_24_15_port, REGISTERS_24_14_port, REGISTERS_24_13_port, 
      REGISTERS_24_12_port, REGISTERS_24_11_port, REGISTERS_24_10_port, 
      REGISTERS_24_9_port, REGISTERS_24_8_port, REGISTERS_24_7_port, 
      REGISTERS_24_6_port, REGISTERS_24_5_port, REGISTERS_24_4_port, 
      REGISTERS_24_3_port, REGISTERS_24_2_port, REGISTERS_24_1_port, 
      REGISTERS_24_0_port, REGISTERS_25_63_port, REGISTERS_25_62_port, 
      REGISTERS_25_61_port, REGISTERS_25_60_port, REGISTERS_25_59_port, 
      REGISTERS_25_58_port, REGISTERS_25_57_port, REGISTERS_25_56_port, 
      REGISTERS_25_55_port, REGISTERS_25_54_port, REGISTERS_25_53_port, 
      REGISTERS_25_52_port, REGISTERS_25_51_port, REGISTERS_25_50_port, 
      REGISTERS_25_49_port, REGISTERS_25_48_port, REGISTERS_25_47_port, 
      REGISTERS_25_46_port, REGISTERS_25_45_port, REGISTERS_25_44_port, 
      REGISTERS_25_43_port, REGISTERS_25_42_port, REGISTERS_25_41_port, 
      REGISTERS_25_40_port, REGISTERS_25_39_port, REGISTERS_25_38_port, 
      REGISTERS_25_37_port, REGISTERS_25_36_port, REGISTERS_25_35_port, 
      REGISTERS_25_34_port, REGISTERS_25_33_port, REGISTERS_25_32_port, 
      REGISTERS_25_31_port, REGISTERS_25_30_port, REGISTERS_25_29_port, 
      REGISTERS_25_28_port, REGISTERS_25_27_port, REGISTERS_25_26_port, 
      REGISTERS_25_25_port, REGISTERS_25_24_port, REGISTERS_25_23_port, 
      REGISTERS_25_22_port, REGISTERS_25_21_port, REGISTERS_25_20_port, 
      REGISTERS_25_19_port, REGISTERS_25_18_port, REGISTERS_25_17_port, 
      REGISTERS_25_16_port, REGISTERS_25_15_port, REGISTERS_25_14_port, 
      REGISTERS_25_13_port, REGISTERS_25_12_port, REGISTERS_25_11_port, 
      REGISTERS_25_10_port, REGISTERS_25_9_port, REGISTERS_25_8_port, 
      REGISTERS_25_7_port, REGISTERS_25_6_port, REGISTERS_25_5_port, 
      REGISTERS_25_4_port, REGISTERS_25_3_port, REGISTERS_25_2_port, 
      REGISTERS_25_1_port, REGISTERS_25_0_port, REGISTERS_26_63_port, 
      REGISTERS_26_62_port, REGISTERS_26_61_port, REGISTERS_26_60_port, 
      REGISTERS_26_59_port, REGISTERS_26_58_port, REGISTERS_26_57_port, 
      REGISTERS_26_56_port, REGISTERS_26_55_port, REGISTERS_26_54_port, 
      REGISTERS_26_53_port, REGISTERS_26_52_port, REGISTERS_26_51_port, 
      REGISTERS_26_50_port, REGISTERS_26_49_port, REGISTERS_26_48_port, 
      REGISTERS_26_47_port, REGISTERS_26_46_port, REGISTERS_26_45_port, 
      REGISTERS_26_44_port, REGISTERS_26_43_port, REGISTERS_26_42_port, 
      REGISTERS_26_41_port, REGISTERS_26_40_port, REGISTERS_26_39_port, 
      REGISTERS_26_38_port, REGISTERS_26_37_port, REGISTERS_26_36_port, 
      REGISTERS_26_35_port, REGISTERS_26_34_port, REGISTERS_26_33_port, 
      REGISTERS_26_32_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_63_port, REGISTERS_27_62_port, REGISTERS_27_61_port, 
      REGISTERS_27_60_port, REGISTERS_27_59_port, REGISTERS_27_58_port, 
      REGISTERS_27_57_port, REGISTERS_27_56_port, REGISTERS_27_55_port, 
      REGISTERS_27_54_port, REGISTERS_27_53_port, REGISTERS_27_52_port, 
      REGISTERS_27_51_port, REGISTERS_27_50_port, REGISTERS_27_49_port, 
      REGISTERS_27_48_port, REGISTERS_27_47_port, REGISTERS_27_46_port, 
      REGISTERS_27_45_port, REGISTERS_27_44_port, REGISTERS_27_43_port, 
      REGISTERS_27_42_port, REGISTERS_27_41_port, REGISTERS_27_40_port, 
      REGISTERS_27_39_port, REGISTERS_27_38_port, REGISTERS_27_37_port, 
      REGISTERS_27_36_port, REGISTERS_27_35_port, REGISTERS_27_34_port, 
      REGISTERS_27_33_port, REGISTERS_27_32_port, REGISTERS_27_31_port, 
      REGISTERS_27_30_port, REGISTERS_27_29_port, REGISTERS_27_28_port, 
      REGISTERS_27_27_port, REGISTERS_27_26_port, REGISTERS_27_25_port, 
      REGISTERS_27_24_port, REGISTERS_27_23_port, REGISTERS_27_22_port, 
      REGISTERS_27_21_port, REGISTERS_27_20_port, REGISTERS_27_19_port, 
      REGISTERS_27_18_port, REGISTERS_27_17_port, REGISTERS_27_16_port, 
      REGISTERS_27_15_port, REGISTERS_27_14_port, REGISTERS_27_13_port, 
      REGISTERS_27_12_port, REGISTERS_27_11_port, REGISTERS_27_10_port, 
      REGISTERS_27_9_port, REGISTERS_27_8_port, REGISTERS_27_7_port, 
      REGISTERS_27_6_port, REGISTERS_27_5_port, REGISTERS_27_4_port, 
      REGISTERS_27_3_port, REGISTERS_27_2_port, REGISTERS_27_1_port, 
      REGISTERS_27_0_port, REGISTERS_28_63_port, REGISTERS_28_62_port, 
      REGISTERS_28_61_port, REGISTERS_28_60_port, REGISTERS_28_59_port, 
      REGISTERS_28_58_port, REGISTERS_28_57_port, REGISTERS_28_56_port, 
      REGISTERS_28_55_port, REGISTERS_28_54_port, REGISTERS_28_53_port, 
      REGISTERS_28_52_port, REGISTERS_28_51_port, REGISTERS_28_50_port, 
      REGISTERS_28_49_port, REGISTERS_28_48_port, REGISTERS_28_47_port, 
      REGISTERS_28_46_port, REGISTERS_28_45_port, REGISTERS_28_44_port, 
      REGISTERS_28_43_port, REGISTERS_28_42_port, REGISTERS_28_41_port, 
      REGISTERS_28_40_port, REGISTERS_28_39_port, REGISTERS_28_38_port, 
      REGISTERS_28_37_port, REGISTERS_28_36_port, REGISTERS_28_35_port, 
      REGISTERS_28_34_port, REGISTERS_28_33_port, REGISTERS_28_32_port, 
      REGISTERS_28_31_port, REGISTERS_28_30_port, REGISTERS_28_29_port, 
      REGISTERS_28_28_port, REGISTERS_28_27_port, REGISTERS_28_26_port, 
      REGISTERS_28_25_port, REGISTERS_28_24_port, REGISTERS_28_23_port, 
      REGISTERS_28_22_port, REGISTERS_28_21_port, REGISTERS_28_20_port, 
      REGISTERS_28_19_port, REGISTERS_28_18_port, REGISTERS_28_17_port, 
      REGISTERS_28_16_port, REGISTERS_28_15_port, REGISTERS_28_14_port, 
      REGISTERS_28_13_port, REGISTERS_28_12_port, REGISTERS_28_11_port, 
      REGISTERS_28_10_port, REGISTERS_28_9_port, REGISTERS_28_8_port, 
      REGISTERS_28_7_port, REGISTERS_28_6_port, REGISTERS_28_5_port, 
      REGISTERS_28_4_port, REGISTERS_28_3_port, REGISTERS_28_2_port, 
      REGISTERS_28_1_port, REGISTERS_28_0_port, REGISTERS_29_63_port, 
      REGISTERS_29_62_port, REGISTERS_29_61_port, REGISTERS_29_60_port, 
      REGISTERS_29_59_port, REGISTERS_29_58_port, REGISTERS_29_57_port, 
      REGISTERS_29_56_port, REGISTERS_29_55_port, REGISTERS_29_54_port, 
      REGISTERS_29_53_port, REGISTERS_29_52_port, REGISTERS_29_51_port, 
      REGISTERS_29_50_port, REGISTERS_29_49_port, REGISTERS_29_48_port, 
      REGISTERS_29_47_port, REGISTERS_29_46_port, REGISTERS_29_45_port, 
      REGISTERS_29_44_port, REGISTERS_29_43_port, REGISTERS_29_42_port, 
      REGISTERS_29_41_port, REGISTERS_29_40_port, REGISTERS_29_39_port, 
      REGISTERS_29_38_port, REGISTERS_29_37_port, REGISTERS_29_36_port, 
      REGISTERS_29_35_port, REGISTERS_29_34_port, REGISTERS_29_33_port, 
      REGISTERS_29_32_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_63_port, REGISTERS_30_62_port, REGISTERS_30_61_port, 
      REGISTERS_30_60_port, REGISTERS_30_59_port, REGISTERS_30_58_port, 
      REGISTERS_30_57_port, REGISTERS_30_56_port, REGISTERS_30_55_port, 
      REGISTERS_30_54_port, REGISTERS_30_53_port, REGISTERS_30_52_port, 
      REGISTERS_30_51_port, REGISTERS_30_50_port, REGISTERS_30_49_port, 
      REGISTERS_30_48_port, REGISTERS_30_47_port, REGISTERS_30_46_port, 
      REGISTERS_30_45_port, REGISTERS_30_44_port, REGISTERS_30_43_port, 
      REGISTERS_30_42_port, REGISTERS_30_41_port, REGISTERS_30_40_port, 
      REGISTERS_30_39_port, REGISTERS_30_38_port, REGISTERS_30_37_port, 
      REGISTERS_30_36_port, REGISTERS_30_35_port, REGISTERS_30_34_port, 
      REGISTERS_30_33_port, REGISTERS_30_32_port, REGISTERS_30_31_port, 
      REGISTERS_30_30_port, REGISTERS_30_29_port, REGISTERS_30_28_port, 
      REGISTERS_30_27_port, REGISTERS_30_26_port, REGISTERS_30_25_port, 
      REGISTERS_30_24_port, REGISTERS_30_23_port, REGISTERS_30_22_port, 
      REGISTERS_30_21_port, REGISTERS_30_20_port, REGISTERS_30_19_port, 
      REGISTERS_30_18_port, REGISTERS_30_17_port, REGISTERS_30_16_port, 
      REGISTERS_30_15_port, REGISTERS_30_14_port, REGISTERS_30_13_port, 
      REGISTERS_30_12_port, REGISTERS_30_11_port, REGISTERS_30_10_port, 
      REGISTERS_30_9_port, REGISTERS_30_8_port, REGISTERS_30_7_port, 
      REGISTERS_30_6_port, REGISTERS_30_5_port, REGISTERS_30_4_port, 
      REGISTERS_30_3_port, REGISTERS_30_2_port, REGISTERS_30_1_port, 
      REGISTERS_30_0_port, REGISTERS_31_63_port, REGISTERS_31_62_port, 
      REGISTERS_31_61_port, REGISTERS_31_60_port, REGISTERS_31_59_port, 
      REGISTERS_31_58_port, REGISTERS_31_57_port, REGISTERS_31_56_port, 
      REGISTERS_31_55_port, REGISTERS_31_54_port, REGISTERS_31_53_port, 
      REGISTERS_31_52_port, REGISTERS_31_51_port, REGISTERS_31_50_port, 
      REGISTERS_31_49_port, REGISTERS_31_48_port, REGISTERS_31_47_port, 
      REGISTERS_31_46_port, REGISTERS_31_45_port, REGISTERS_31_44_port, 
      REGISTERS_31_43_port, REGISTERS_31_42_port, REGISTERS_31_41_port, 
      REGISTERS_31_40_port, REGISTERS_31_39_port, REGISTERS_31_38_port, 
      REGISTERS_31_37_port, REGISTERS_31_36_port, REGISTERS_31_35_port, 
      REGISTERS_31_34_port, REGISTERS_31_33_port, REGISTERS_31_32_port, 
      REGISTERS_31_31_port, REGISTERS_31_30_port, REGISTERS_31_29_port, 
      REGISTERS_31_28_port, REGISTERS_31_27_port, REGISTERS_31_26_port, 
      REGISTERS_31_25_port, REGISTERS_31_24_port, REGISTERS_31_23_port, 
      REGISTERS_31_22_port, REGISTERS_31_21_port, REGISTERS_31_20_port, 
      REGISTERS_31_19_port, REGISTERS_31_18_port, REGISTERS_31_17_port, 
      REGISTERS_31_16_port, REGISTERS_31_15_port, REGISTERS_31_14_port, 
      REGISTERS_31_13_port, REGISTERS_31_12_port, REGISTERS_31_11_port, 
      REGISTERS_31_10_port, REGISTERS_31_9_port, REGISTERS_31_8_port, 
      REGISTERS_31_7_port, REGISTERS_31_6_port, REGISTERS_31_5_port, 
      REGISTERS_31_4_port, REGISTERS_31_3_port, REGISTERS_31_2_port, 
      REGISTERS_31_1_port, REGISTERS_31_0_port, N96, N97, N98, N99, N100, N101,
      N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, 
      N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, 
      N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, 
      N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, 
      N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N225, N226, 
      N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, 
      N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, 
      N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, 
      N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, 
      N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, 
      N287, N288, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464
      , n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, 
      n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, 
      n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, 
      n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, 
      n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, 
      n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, 
      n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, 
      n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, 
      n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, 
      n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, 
      n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, 
      n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, 
      n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, 
      n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, 
      n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, 
      n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, 
      n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, 
      n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, 
      n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, 
      n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, 
      n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, 
      n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, 
      n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, 
      n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, 
      n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, 
      n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, 
      n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, 
      n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, 
      n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, 
      n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, 
      n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, 
      n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, 
      n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, 
      n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, 
      n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, 
      n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, 
      n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, 
      n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, 
      n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, 
      n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, 
      n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, 
      n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, 
      n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, 
      n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, 
      n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, 
      n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, 
      n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, 
      n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, 
      n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, 
      n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, 
      n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, 
      n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, 
      n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, 
      n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, 
      n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, 
      n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, 
      n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, 
      n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, 
      n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, 
      n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, 
      n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, 
      n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, 
      n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, 
      n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, 
      n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, 
      n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, 
      n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, 
      n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, 
      n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, 
      n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, 
      n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, 
      n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, 
      n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, 
      n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, 
      n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, 
      n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, 
      n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, 
      n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, 
      n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, 
      n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, 
      n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, 
      n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, 
      n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, 
      n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, 
      n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, 
      n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, 
      n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, 
      n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, 
      n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, 
      n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, 
      n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, 
      n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, 
      n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, 
      n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, 
      n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, 
      n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, 
      n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, 
      n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, 
      n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, 
      n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, 
      n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, 
      n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, 
      n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, 
      n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, 
      n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, 
      n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, 
      n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, 
      n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, 
      n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, 
      n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, 
      n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, 
      n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, 
      n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, 
      n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, 
      n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, 
      n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, 
      n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, 
      n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, 
      n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, 
      n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, 
      n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, 
      n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, 
      n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, 
      n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, 
      n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, 
      n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, 
      n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, 
      n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, 
      n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, 
      n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, 
      n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, 
      n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, 
      n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, 
      n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, 
      n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, 
      n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, 
      n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, 
      n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, 
      n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, 
      n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, 
      n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, 
      n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, 
      n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, 
      n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, 
      n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, 
      n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, 
      n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, 
      n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, 
      n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, 
      n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, 
      n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, 
      n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, 
      n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, 
      n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, 
      n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, 
      n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, 
      n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, 
      n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, 
      n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, 
      n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, 
      n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, 
      n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, 
      n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, 
      n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, 
      n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, 
      n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, 
      n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, 
      n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, 
      n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, 
      n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, 
      n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, 
      n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, 
      n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, 
      n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, 
      n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, 
      n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, 
      n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, 
      n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, 
      n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, 
      n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, 
      n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, 
      n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, 
      n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, 
      n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, 
      n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, 
      n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, 
      n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, 
      n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, 
      n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, 
      n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, 
      n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, 
      n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, 
      n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, 
      n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, 
      n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, 
      n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, 
      n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, 
      n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, 
      n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, 
      n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, 
      n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, 
      n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, 
      n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, 
      n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n1, n2, n3
      , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91
      , n92, n93, n94, n95, n96_port, n97_port, n98_port, n99_port, n100_port, 
      n101_port, n102_port, n103_port, n104_port, n105_port, n106_port, 
      n107_port, n108_port, n109_port, n110_port, n111_port, n112_port, 
      n113_port, n114_port, n115_port, n116_port, n117_port, n118_port, 
      n119_port, n120_port, n121_port, n122_port, n123_port, n124_port, 
      n125_port, n126_port, n127_port, n128_port, n129_port, n130_port, 
      n131_port, n132_port, n133_port, n134_port, n135_port, n136_port, 
      n137_port, n138_port, n139_port, n140_port, n141_port, n142_port, 
      n143_port, n144_port, n145_port, n146_port, n147_port, n148_port, 
      n149_port, n150_port, n151_port, n152_port, n153_port, n154_port, 
      n155_port, n156_port, n157_port, n158_port, n159_port, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225_port, n226_port, n227_port, n228_port, n229_port, 
      n230_port, n231_port, n232_port, n233_port, n234_port, n235_port, 
      n236_port, n237_port, n238_port, n239_port, n240_port, n241_port, 
      n242_port, n243_port, n244_port, n245_port, n246_port, n247_port, 
      n248_port, n249_port, n250_port, n251_port, n252_port, n253_port, 
      n254_port, n255_port, n256_port, n257_port, n258_port, n259_port, 
      n260_port, n261_port, n262_port, n263_port, n264_port, n265_port, 
      n266_port, n267_port, n268_port, n269_port, n270_port, n271_port, 
      n272_port, n273_port, n274_port, n275_port, n276_port, n277_port, 
      n278_port, n279_port, n280_port, n281_port, n282_port, n283_port, 
      n284_port, n285_port, n286_port, n287_port, n288_port, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, 
      n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, 
      n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
      n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
      n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
      n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, 
      n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, 
      n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
      n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
      n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, 
      n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
      n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, 
      n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, 
      n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, 
      n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, 
      n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, 
      n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, 
      n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, 
      n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
      n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
      n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
      n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
      n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
      n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
      n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
      n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, 
      n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
      n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, 
      n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
      n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, 
      n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
      n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
      n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, 
      n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, 
      n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, 
      n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, 
      n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, 
      n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, 
      n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
      n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, 
      n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
      n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, 
      n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
      n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, 
      n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
      n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, 
      n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
      n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
      n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, 
      n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, 
      n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, 
      n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, 
      n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, 
      n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, 
      n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, 
      n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
      n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
      n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, 
      n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
      n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
      n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, 
      n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, 
      n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, 
      n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, 
      n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, 
      n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, 
      n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
      n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, 
      n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, 
      n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, 
      n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, 
      n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, 
      n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, 
      n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, 
      n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, 
      n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, 
      n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, 
      n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, 
      n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, 
      n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
      n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, 
      n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, 
      n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, 
      n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, 
      n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, 
      n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, 
      n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
      n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, 
      n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, 
      n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, 
      n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, 
      n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, 
      n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, 
      n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, 
      n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, 
      n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, 
      n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
      n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
      n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
      n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
      n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, 
      n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, 
      n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, 
      n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, 
      n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, 
      n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, 
      n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, 
      n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, 
      n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, 
      n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, 
      n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, 
      n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, 
      n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, 
      n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, 
      n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, 
      n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, 
      n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, 
      n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, 
      n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, 
      n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, 
      n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, 
      n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, 
      n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, 
      n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, 
      n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, 
      n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, 
      n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, 
      n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, 
      n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, 
      n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, 
      n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, 
      n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, 
      n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, 
      n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, 
      n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, 
      n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, 
      n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, 
      n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, 
      n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, 
      n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, 
      n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, 
      n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, 
      n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, 
      n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, 
      n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, 
      n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, 
      n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, 
      n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, 
      n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, 
      n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, 
      n2450, n2451, n2452, n2453, n2454, n2455, n4504, n4505, n4506, n4507, 
      n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, 
      n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, 
      n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, 
      n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, 
      n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, 
      n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, 
      n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, 
      n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, 
      n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, 
      n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, 
      n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, 
      n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, 
      n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, 
      n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, 
      n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, 
      n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, 
      n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, 
      n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, 
      n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, 
      n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, 
      n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, 
      n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, 
      n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, 
      n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, 
      n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, 
      n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, 
      n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, 
      n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, 
      n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, 
      n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, 
      n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, 
      n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, 
      n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, 
      n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, 
      n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, 
      n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, 
      n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, 
      n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, 
      n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, 
      n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, 
      n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, 
      n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, 
      n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, 
      n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, 
      n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, 
      n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, 
      n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, 
      n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, 
      n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, 
      n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, 
      n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, 
      n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, 
      n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, 
      n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, 
      n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, 
      n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, 
      n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, 
      n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, 
      n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, 
      n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, 
      n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, 
      n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, 
      n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, 
      n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, 
      n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, 
      n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, 
      n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, 
      n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, 
      n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, 
      n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, 
      n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, 
      n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, 
      n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, 
      n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, 
      n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, 
      n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, 
      n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, 
      n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, 
      n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, 
      n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, 
      n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, 
      n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, 
      n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, 
      n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, 
      n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, 
      n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, 
      n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, 
      n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, 
      n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, 
      n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, 
      n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, 
      n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, 
      n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, 
      n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, 
      n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, 
      n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, 
      n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, 
      n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, 
      n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, 
      n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, 
      n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, 
      n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, 
      n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, 
      n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, 
      n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, 
      n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, 
      n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, 
      n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, 
      n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, 
      n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, 
      n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, 
      n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, 
      n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, 
      n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, 
      n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, 
      n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, 
      n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, 
      n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, 
      n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, 
      n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, 
      n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, 
      n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, 
      n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, 
      n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, 
      n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, 
      n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, 
      n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, 
      n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, 
      n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, 
      n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, 
      n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, 
      n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, 
      n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, 
      n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, 
      n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, 
      n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, 
      n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, 
      n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, 
      n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, 
      n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, 
      n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, 
      n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, 
      n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, 
      n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, 
      n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, 
      n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, 
      n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, 
      n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, 
      n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, 
      n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, 
      n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, 
      n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, 
      n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, 
      n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, 
      n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, 
      n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, 
      n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, 
      n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, 
      n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, 
      n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, 
      n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, 
      n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, 
      n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, 
      n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, 
      n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, 
      n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, 
      n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, 
      n6178, n6179, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, 
      n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, 
      n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, 
      n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, 
      n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, 
      n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, 
      n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, 
      n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, 
      n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, 
      n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, 
      n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, 
      n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, 
      n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, 
      n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, 
      n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, 
      n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, 
      n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, 
      n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, 
      n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, 
      n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, 
      n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, 
      n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, 
      n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, 
      n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, 
      n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, 
      n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, 
      n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, 
      n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, 
      n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, 
      n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, 
      n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, 
      n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, 
      n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, 
      n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, 
      n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, 
      n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, 
      n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, 
      n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, 
      n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, 
      n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, 
      n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, 
      n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, 
      n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, 
      n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, 
      n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, 
      n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, 
      n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, 
      n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, 
      n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, 
      n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, 
      n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, 
      n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, 
      n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, 
      n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, 
      n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, 
      n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, 
      n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, 
      n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, 
      n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, 
      n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, 
      n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, 
      n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, 
      n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, 
      n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, 
      n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, 
      n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, 
      n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, 
      n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, 
      n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, 
      n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, 
      n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, 
      n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, 
      n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, 
      n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, 
      n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, 
      n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, 
      n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, 
      n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, 
      n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, 
      n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, 
      n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, 
      n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, 
      n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, 
      n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, 
      n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, 
      n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, 
      n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, 
      n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, 
      n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, 
      n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, 
      n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, 
      n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, 
      n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, 
      n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, 
      n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, 
      n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, 
      n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, 
      n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, 
      n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, 
      n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, 
      n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, 
      n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, 
      n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, 
      n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, 
      n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, 
      n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, 
      n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, 
      n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, 
      n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, 
      n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, 
      n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, 
      n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, 
      n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, 
      n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, 
      n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, 
      n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, 
      n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, 
      n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, 
      n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, 
      n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, 
      n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, 
      n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, 
      n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, 
      n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, 
      n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, 
      n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, 
      n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, 
      n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, 
      n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, 
      n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, 
      n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, 
      n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, 
      n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, 
      n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, 
      n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, 
      n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, 
      n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, 
      n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, 
      n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, 
      n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, 
      n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, 
      n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, 
      n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, 
      n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, 
      n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, 
      n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, 
      n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, 
      n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, 
      n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, 
      n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, 
      n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, 
      n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, 
      n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, 
      n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, 
      n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, 
      n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, 
      n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, 
      n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, 
      n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, 
      n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, 
      n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, 
      n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, 
      n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, 
      n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, 
      n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, 
      n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, n_3051 : std_logic;

begin
   
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n4503, CK => n804, Q => 
                           REGISTERS_0_63_port, QN => n_1004);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n4502, CK => n804, Q => 
                           REGISTERS_0_62_port, QN => n_1005);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n4501, CK => n804, Q => 
                           REGISTERS_0_61_port, QN => n_1006);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n4500, CK => n805, Q => 
                           REGISTERS_0_60_port, QN => n_1007);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n4499, CK => n805, Q => 
                           REGISTERS_0_59_port, QN => n_1008);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n4498, CK => n805, Q => 
                           REGISTERS_0_58_port, QN => n_1009);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n4497, CK => n805, Q => 
                           REGISTERS_0_57_port, QN => n_1010);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n4496, CK => n805, Q => 
                           REGISTERS_0_56_port, QN => n_1011);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n4495, CK => n805, Q => 
                           REGISTERS_0_55_port, QN => n_1012);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n4494, CK => n805, Q => 
                           REGISTERS_0_54_port, QN => n_1013);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n4493, CK => n805, Q => 
                           REGISTERS_0_53_port, QN => n_1014);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n4492, CK => n805, Q => 
                           REGISTERS_0_52_port, QN => n_1015);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n4491, CK => n805, Q => 
                           REGISTERS_0_51_port, QN => n_1016);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n4490, CK => n805, Q => 
                           REGISTERS_0_50_port, QN => n_1017);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n4489, CK => n806, Q => 
                           REGISTERS_0_49_port, QN => n_1018);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n4488, CK => n806, Q => 
                           REGISTERS_0_48_port, QN => n_1019);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n4487, CK => n806, Q => 
                           REGISTERS_0_47_port, QN => n_1020);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n4486, CK => n806, Q => 
                           REGISTERS_0_46_port, QN => n_1021);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n4485, CK => n806, Q => 
                           REGISTERS_0_45_port, QN => n_1022);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n4484, CK => n806, Q => 
                           REGISTERS_0_44_port, QN => n_1023);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n4483, CK => n806, Q => 
                           REGISTERS_0_43_port, QN => n_1024);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n4482, CK => n806, Q => 
                           REGISTERS_0_42_port, QN => n_1025);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n4481, CK => n806, Q => 
                           REGISTERS_0_41_port, QN => n_1026);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n4480, CK => n806, Q => 
                           REGISTERS_0_40_port, QN => n_1027);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n4479, CK => n806, Q => 
                           REGISTERS_0_39_port, QN => n_1028);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n4478, CK => n807, Q => 
                           REGISTERS_0_38_port, QN => n_1029);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n4477, CK => n807, Q => 
                           REGISTERS_0_37_port, QN => n_1030);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n4476, CK => n807, Q => 
                           REGISTERS_0_36_port, QN => n_1031);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n4475, CK => n807, Q => 
                           REGISTERS_0_35_port, QN => n_1032);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n4474, CK => n807, Q => 
                           REGISTERS_0_34_port, QN => n_1033);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n4473, CK => n807, Q => 
                           REGISTERS_0_33_port, QN => n_1034);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n4472, CK => n807, Q => 
                           REGISTERS_0_32_port, QN => n_1035);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n4471, CK => n807, Q => 
                           REGISTERS_0_31_port, QN => n_1036);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n4470, CK => n807, Q => 
                           REGISTERS_0_30_port, QN => n_1037);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n4469, CK => n807, Q => 
                           REGISTERS_0_29_port, QN => n_1038);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n4468, CK => n807, Q => 
                           REGISTERS_0_28_port, QN => n_1039);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n4467, CK => n808, Q => 
                           REGISTERS_0_27_port, QN => n_1040);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n4466, CK => n808, Q => 
                           REGISTERS_0_26_port, QN => n_1041);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n4465, CK => n808, Q => 
                           REGISTERS_0_25_port, QN => n_1042);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n4464, CK => n808, Q => 
                           REGISTERS_0_24_port, QN => n_1043);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n4463, CK => n808, Q => 
                           REGISTERS_0_23_port, QN => n_1044);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n4462, CK => n808, Q => 
                           REGISTERS_0_22_port, QN => n_1045);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n4461, CK => n808, Q => 
                           REGISTERS_0_21_port, QN => n_1046);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n4460, CK => n808, Q => 
                           REGISTERS_0_20_port, QN => n_1047);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n4459, CK => n808, Q => 
                           REGISTERS_0_19_port, QN => n_1048);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n4458, CK => n808, Q => 
                           REGISTERS_0_18_port, QN => n_1049);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n4457, CK => n808, Q => 
                           REGISTERS_0_17_port, QN => n_1050);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n4456, CK => n809, Q => 
                           REGISTERS_0_16_port, QN => n_1051);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n4455, CK => n809, Q => 
                           REGISTERS_0_15_port, QN => n_1052);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n4454, CK => n809, Q => 
                           REGISTERS_0_14_port, QN => n_1053);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n4453, CK => n809, Q => 
                           REGISTERS_0_13_port, QN => n_1054);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n4452, CK => n809, Q => 
                           REGISTERS_0_12_port, QN => n_1055);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n4451, CK => n809, Q => 
                           REGISTERS_0_11_port, QN => n_1056);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n4450, CK => n809, Q => 
                           REGISTERS_0_10_port, QN => n_1057);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n4449, CK => n809, Q => 
                           REGISTERS_0_9_port, QN => n_1058);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n4448, CK => n809, Q => 
                           REGISTERS_0_8_port, QN => n_1059);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n4447, CK => n809, Q => 
                           REGISTERS_0_7_port, QN => n_1060);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n4446, CK => n809, Q => 
                           REGISTERS_0_6_port, QN => n_1061);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n4445, CK => n810, Q => 
                           REGISTERS_0_5_port, QN => n_1062);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n4444, CK => n810, Q => 
                           REGISTERS_0_4_port, QN => n_1063);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n4443, CK => n810, Q => 
                           REGISTERS_0_3_port, QN => n_1064);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n4442, CK => n810, Q => 
                           REGISTERS_0_2_port, QN => n_1065);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n4441, CK => n810, Q => 
                           REGISTERS_0_1_port, QN => n_1066);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n4440, CK => n810, Q => 
                           REGISTERS_0_0_port, QN => n_1067);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n4439, CK => n810, Q => 
                           REGISTERS_1_63_port, QN => n_1068);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n4438, CK => n810, Q => 
                           REGISTERS_1_62_port, QN => n_1069);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n4437, CK => n810, Q => 
                           REGISTERS_1_61_port, QN => n_1070);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n4436, CK => n810, Q => 
                           REGISTERS_1_60_port, QN => n_1071);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n4435, CK => n810, Q => 
                           REGISTERS_1_59_port, QN => n_1072);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n4434, CK => n811, Q => 
                           REGISTERS_1_58_port, QN => n_1073);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n4433, CK => n811, Q => 
                           REGISTERS_1_57_port, QN => n_1074);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n4432, CK => n811, Q => 
                           REGISTERS_1_56_port, QN => n_1075);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n4431, CK => n811, Q => 
                           REGISTERS_1_55_port, QN => n_1076);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n4430, CK => n811, Q => 
                           REGISTERS_1_54_port, QN => n_1077);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n4429, CK => n811, Q => 
                           REGISTERS_1_53_port, QN => n_1078);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n4428, CK => n811, Q => 
                           REGISTERS_1_52_port, QN => n_1079);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n4427, CK => n811, Q => 
                           REGISTERS_1_51_port, QN => n_1080);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n4426, CK => n811, Q => 
                           REGISTERS_1_50_port, QN => n_1081);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n4425, CK => n811, Q => 
                           REGISTERS_1_49_port, QN => n_1082);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n4424, CK => n811, Q => 
                           REGISTERS_1_48_port, QN => n_1083);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n4423, CK => n812, Q => 
                           REGISTERS_1_47_port, QN => n_1084);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n4422, CK => n812, Q => 
                           REGISTERS_1_46_port, QN => n_1085);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n4421, CK => n812, Q => 
                           REGISTERS_1_45_port, QN => n_1086);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n4420, CK => n812, Q => 
                           REGISTERS_1_44_port, QN => n_1087);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n4419, CK => n812, Q => 
                           REGISTERS_1_43_port, QN => n_1088);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n4418, CK => n812, Q => 
                           REGISTERS_1_42_port, QN => n_1089);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n4417, CK => n812, Q => 
                           REGISTERS_1_41_port, QN => n_1090);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n4416, CK => n812, Q => 
                           REGISTERS_1_40_port, QN => n_1091);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n4415, CK => n812, Q => 
                           REGISTERS_1_39_port, QN => n_1092);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n4414, CK => n812, Q => 
                           REGISTERS_1_38_port, QN => n_1093);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n4413, CK => n812, Q => 
                           REGISTERS_1_37_port, QN => n_1094);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n4412, CK => n813, Q => 
                           REGISTERS_1_36_port, QN => n_1095);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n4411, CK => n813, Q => 
                           REGISTERS_1_35_port, QN => n_1096);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n4410, CK => n813, Q => 
                           REGISTERS_1_34_port, QN => n_1097);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n4409, CK => n813, Q => 
                           REGISTERS_1_33_port, QN => n_1098);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n4408, CK => n813, Q => 
                           REGISTERS_1_32_port, QN => n_1099);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n4407, CK => n813, Q => 
                           REGISTERS_1_31_port, QN => n_1100);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n4406, CK => n813, Q => 
                           REGISTERS_1_30_port, QN => n_1101);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n4405, CK => n813, Q => 
                           REGISTERS_1_29_port, QN => n_1102);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n4404, CK => n813, Q => 
                           REGISTERS_1_28_port, QN => n_1103);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n4403, CK => n813, Q => 
                           REGISTERS_1_27_port, QN => n_1104);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n4402, CK => n813, Q => 
                           REGISTERS_1_26_port, QN => n_1105);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n4401, CK => n814, Q => 
                           REGISTERS_1_25_port, QN => n_1106);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n4400, CK => n814, Q => 
                           REGISTERS_1_24_port, QN => n_1107);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n4399, CK => n814, Q => 
                           REGISTERS_1_23_port, QN => n_1108);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n4398, CK => n814, Q => 
                           REGISTERS_1_22_port, QN => n_1109);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n4397, CK => n814, Q => 
                           REGISTERS_1_21_port, QN => n_1110);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n4396, CK => n814, Q => 
                           REGISTERS_1_20_port, QN => n_1111);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n4395, CK => n814, Q => 
                           REGISTERS_1_19_port, QN => n_1112);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n4394, CK => n814, Q => 
                           REGISTERS_1_18_port, QN => n_1113);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n4393, CK => n814, Q => 
                           REGISTERS_1_17_port, QN => n_1114);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n4392, CK => n814, Q => 
                           REGISTERS_1_16_port, QN => n_1115);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n4391, CK => n814, Q => 
                           REGISTERS_1_15_port, QN => n_1116);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n4390, CK => n815, Q => 
                           REGISTERS_1_14_port, QN => n_1117);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n4389, CK => n815, Q => 
                           REGISTERS_1_13_port, QN => n_1118);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n4388, CK => n815, Q => 
                           REGISTERS_1_12_port, QN => n_1119);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n4387, CK => n815, Q => 
                           REGISTERS_1_11_port, QN => n_1120);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n4386, CK => n815, Q => 
                           REGISTERS_1_10_port, QN => n_1121);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n4385, CK => n815, Q => 
                           REGISTERS_1_9_port, QN => n_1122);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n4384, CK => n815, Q => 
                           REGISTERS_1_8_port, QN => n_1123);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n4383, CK => n815, Q => 
                           REGISTERS_1_7_port, QN => n_1124);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n4382, CK => n815, Q => 
                           REGISTERS_1_6_port, QN => n_1125);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n4381, CK => n815, Q => 
                           REGISTERS_1_5_port, QN => n_1126);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n4380, CK => n815, Q => 
                           REGISTERS_1_4_port, QN => n_1127);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n4379, CK => n816, Q => 
                           REGISTERS_1_3_port, QN => n_1128);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n4378, CK => n816, Q => 
                           REGISTERS_1_2_port, QN => n_1129);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n4377, CK => n816, Q => 
                           REGISTERS_1_1_port, QN => n_1130);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n4376, CK => n816, Q => 
                           REGISTERS_1_0_port, QN => n_1131);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n4375, CK => n816, Q => 
                           REGISTERS_2_63_port, QN => n_1132);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n4374, CK => n816, Q => 
                           REGISTERS_2_62_port, QN => n_1133);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n4373, CK => n816, Q => 
                           REGISTERS_2_61_port, QN => n_1134);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n4372, CK => n816, Q => 
                           REGISTERS_2_60_port, QN => n_1135);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n4371, CK => n816, Q => 
                           REGISTERS_2_59_port, QN => n_1136);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n4370, CK => n816, Q => 
                           REGISTERS_2_58_port, QN => n_1137);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n4369, CK => n816, Q => 
                           REGISTERS_2_57_port, QN => n_1138);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n4368, CK => n817, Q => 
                           REGISTERS_2_56_port, QN => n_1139);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n4367, CK => n817, Q => 
                           REGISTERS_2_55_port, QN => n_1140);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n4366, CK => n817, Q => 
                           REGISTERS_2_54_port, QN => n_1141);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n4365, CK => n817, Q => 
                           REGISTERS_2_53_port, QN => n_1142);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n4364, CK => n817, Q => 
                           REGISTERS_2_52_port, QN => n_1143);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n4363, CK => n817, Q => 
                           REGISTERS_2_51_port, QN => n_1144);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n4362, CK => n817, Q => 
                           REGISTERS_2_50_port, QN => n_1145);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n4361, CK => n817, Q => 
                           REGISTERS_2_49_port, QN => n_1146);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n4360, CK => n817, Q => 
                           REGISTERS_2_48_port, QN => n_1147);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n4359, CK => n817, Q => 
                           REGISTERS_2_47_port, QN => n_1148);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n4358, CK => n817, Q => 
                           REGISTERS_2_46_port, QN => n_1149);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n4357, CK => n818, Q => 
                           REGISTERS_2_45_port, QN => n_1150);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n4356, CK => n818, Q => 
                           REGISTERS_2_44_port, QN => n_1151);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n4355, CK => n818, Q => 
                           REGISTERS_2_43_port, QN => n_1152);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n4354, CK => n818, Q => 
                           REGISTERS_2_42_port, QN => n_1153);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n4353, CK => n818, Q => 
                           REGISTERS_2_41_port, QN => n_1154);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n4352, CK => n818, Q => 
                           REGISTERS_2_40_port, QN => n_1155);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n4351, CK => n818, Q => 
                           REGISTERS_2_39_port, QN => n_1156);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n4350, CK => n818, Q => 
                           REGISTERS_2_38_port, QN => n_1157);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n4349, CK => n818, Q => 
                           REGISTERS_2_37_port, QN => n_1158);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n4348, CK => n818, Q => 
                           REGISTERS_2_36_port, QN => n_1159);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n4347, CK => n818, Q => 
                           REGISTERS_2_35_port, QN => n_1160);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n4346, CK => n819, Q => 
                           REGISTERS_2_34_port, QN => n_1161);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n4345, CK => n819, Q => 
                           REGISTERS_2_33_port, QN => n_1162);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n4344, CK => n819, Q => 
                           REGISTERS_2_32_port, QN => n_1163);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n4343, CK => n819, Q => 
                           REGISTERS_2_31_port, QN => n_1164);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n4342, CK => n819, Q => 
                           REGISTERS_2_30_port, QN => n_1165);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n4341, CK => n819, Q => 
                           REGISTERS_2_29_port, QN => n_1166);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n4340, CK => n819, Q => 
                           REGISTERS_2_28_port, QN => n_1167);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n4339, CK => n819, Q => 
                           REGISTERS_2_27_port, QN => n_1168);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n4338, CK => n819, Q => 
                           REGISTERS_2_26_port, QN => n_1169);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n4337, CK => n819, Q => 
                           REGISTERS_2_25_port, QN => n_1170);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n4336, CK => n819, Q => 
                           REGISTERS_2_24_port, QN => n_1171);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n4335, CK => n820, Q => 
                           REGISTERS_2_23_port, QN => n_1172);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n4334, CK => n820, Q => 
                           REGISTERS_2_22_port, QN => n_1173);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n4333, CK => n820, Q => 
                           REGISTERS_2_21_port, QN => n_1174);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n4332, CK => n820, Q => 
                           REGISTERS_2_20_port, QN => n_1175);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n4331, CK => n820, Q => 
                           REGISTERS_2_19_port, QN => n_1176);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n4330, CK => n820, Q => 
                           REGISTERS_2_18_port, QN => n_1177);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n4329, CK => n820, Q => 
                           REGISTERS_2_17_port, QN => n_1178);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n4328, CK => n820, Q => 
                           REGISTERS_2_16_port, QN => n_1179);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n4327, CK => n820, Q => 
                           REGISTERS_2_15_port, QN => n_1180);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n4326, CK => n820, Q => 
                           REGISTERS_2_14_port, QN => n_1181);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n4325, CK => n820, Q => 
                           REGISTERS_2_13_port, QN => n_1182);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n4324, CK => n821, Q => 
                           REGISTERS_2_12_port, QN => n_1183);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n4323, CK => n821, Q => 
                           REGISTERS_2_11_port, QN => n_1184);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n4322, CK => n821, Q => 
                           REGISTERS_2_10_port, QN => n_1185);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n4321, CK => n821, Q => 
                           REGISTERS_2_9_port, QN => n_1186);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n4320, CK => n821, Q => 
                           REGISTERS_2_8_port, QN => n_1187);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n4319, CK => n821, Q => 
                           REGISTERS_2_7_port, QN => n_1188);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n4318, CK => n821, Q => 
                           REGISTERS_2_6_port, QN => n_1189);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n4317, CK => n821, Q => 
                           REGISTERS_2_5_port, QN => n_1190);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n4316, CK => n821, Q => 
                           REGISTERS_2_4_port, QN => n_1191);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n4315, CK => n821, Q => 
                           REGISTERS_2_3_port, QN => n_1192);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n4314, CK => n821, Q => 
                           REGISTERS_2_2_port, QN => n_1193);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n4313, CK => n822, Q => 
                           REGISTERS_2_1_port, QN => n_1194);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n4312, CK => n822, Q => 
                           REGISTERS_2_0_port, QN => n_1195);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n4311, CK => n822, Q => 
                           REGISTERS_3_63_port, QN => n_1196);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n4310, CK => n822, Q => 
                           REGISTERS_3_62_port, QN => n_1197);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n4309, CK => n822, Q => 
                           REGISTERS_3_61_port, QN => n_1198);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n4308, CK => n822, Q => 
                           REGISTERS_3_60_port, QN => n_1199);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n4307, CK => n822, Q => 
                           REGISTERS_3_59_port, QN => n_1200);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n4306, CK => n822, Q => 
                           REGISTERS_3_58_port, QN => n_1201);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n4305, CK => n822, Q => 
                           REGISTERS_3_57_port, QN => n_1202);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n4304, CK => n822, Q => 
                           REGISTERS_3_56_port, QN => n_1203);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n4303, CK => n822, Q => 
                           REGISTERS_3_55_port, QN => n_1204);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n4302, CK => n823, Q => 
                           REGISTERS_3_54_port, QN => n_1205);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n4301, CK => n823, Q => 
                           REGISTERS_3_53_port, QN => n_1206);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n4300, CK => n823, Q => 
                           REGISTERS_3_52_port, QN => n_1207);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n4299, CK => n823, Q => 
                           REGISTERS_3_51_port, QN => n_1208);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n4298, CK => n823, Q => 
                           REGISTERS_3_50_port, QN => n_1209);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n4297, CK => n823, Q => 
                           REGISTERS_3_49_port, QN => n_1210);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n4296, CK => n823, Q => 
                           REGISTERS_3_48_port, QN => n_1211);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n4295, CK => n823, Q => 
                           REGISTERS_3_47_port, QN => n_1212);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n4294, CK => n823, Q => 
                           REGISTERS_3_46_port, QN => n_1213);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n4293, CK => n823, Q => 
                           REGISTERS_3_45_port, QN => n_1214);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n4292, CK => n823, Q => 
                           REGISTERS_3_44_port, QN => n_1215);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n4291, CK => n824, Q => 
                           REGISTERS_3_43_port, QN => n_1216);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n4290, CK => n824, Q => 
                           REGISTERS_3_42_port, QN => n_1217);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n4289, CK => n824, Q => 
                           REGISTERS_3_41_port, QN => n_1218);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n4288, CK => n824, Q => 
                           REGISTERS_3_40_port, QN => n_1219);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n4287, CK => n824, Q => 
                           REGISTERS_3_39_port, QN => n_1220);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n4286, CK => n824, Q => 
                           REGISTERS_3_38_port, QN => n_1221);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n4285, CK => n824, Q => 
                           REGISTERS_3_37_port, QN => n_1222);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n4284, CK => n824, Q => 
                           REGISTERS_3_36_port, QN => n_1223);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n4283, CK => n824, Q => 
                           REGISTERS_3_35_port, QN => n_1224);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n4282, CK => n824, Q => 
                           REGISTERS_3_34_port, QN => n_1225);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n4281, CK => n824, Q => 
                           REGISTERS_3_33_port, QN => n_1226);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n4280, CK => n825, Q => 
                           REGISTERS_3_32_port, QN => n_1227);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n4279, CK => n825, Q => 
                           REGISTERS_3_31_port, QN => n_1228);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n4278, CK => n825, Q => 
                           REGISTERS_3_30_port, QN => n_1229);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n4277, CK => n825, Q => 
                           REGISTERS_3_29_port, QN => n_1230);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n4276, CK => n825, Q => 
                           REGISTERS_3_28_port, QN => n_1231);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n4275, CK => n825, Q => 
                           REGISTERS_3_27_port, QN => n_1232);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n4274, CK => n825, Q => 
                           REGISTERS_3_26_port, QN => n_1233);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n4273, CK => n825, Q => 
                           REGISTERS_3_25_port, QN => n_1234);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n4272, CK => n825, Q => 
                           REGISTERS_3_24_port, QN => n_1235);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n4271, CK => n825, Q => 
                           REGISTERS_3_23_port, QN => n_1236);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n4270, CK => n825, Q => 
                           REGISTERS_3_22_port, QN => n_1237);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n4269, CK => n826, Q => 
                           REGISTERS_3_21_port, QN => n_1238);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n4268, CK => n826, Q => 
                           REGISTERS_3_20_port, QN => n_1239);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n4267, CK => n826, Q => 
                           REGISTERS_3_19_port, QN => n_1240);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n4266, CK => n826, Q => 
                           REGISTERS_3_18_port, QN => n_1241);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n4265, CK => n826, Q => 
                           REGISTERS_3_17_port, QN => n_1242);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n4264, CK => n826, Q => 
                           REGISTERS_3_16_port, QN => n_1243);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n4263, CK => n826, Q => 
                           REGISTERS_3_15_port, QN => n_1244);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n4262, CK => n826, Q => 
                           REGISTERS_3_14_port, QN => n_1245);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n4261, CK => n826, Q => 
                           REGISTERS_3_13_port, QN => n_1246);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n4260, CK => n826, Q => 
                           REGISTERS_3_12_port, QN => n_1247);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n4259, CK => n826, Q => 
                           REGISTERS_3_11_port, QN => n_1248);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n4258, CK => n827, Q => 
                           REGISTERS_3_10_port, QN => n_1249);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n4257, CK => n827, Q => 
                           REGISTERS_3_9_port, QN => n_1250);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n4256, CK => n827, Q => 
                           REGISTERS_3_8_port, QN => n_1251);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n4255, CK => n827, Q => 
                           REGISTERS_3_7_port, QN => n_1252);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n4254, CK => n827, Q => 
                           REGISTERS_3_6_port, QN => n_1253);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n4253, CK => n827, Q => 
                           REGISTERS_3_5_port, QN => n_1254);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n4252, CK => n827, Q => 
                           REGISTERS_3_4_port, QN => n_1255);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n4251, CK => n827, Q => 
                           REGISTERS_3_3_port, QN => n_1256);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n4250, CK => n827, Q => 
                           REGISTERS_3_2_port, QN => n_1257);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n4249, CK => n827, Q => 
                           REGISTERS_3_1_port, QN => n_1258);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n4248, CK => n827, Q => 
                           REGISTERS_3_0_port, QN => n_1259);
   REGISTERS_reg_4_63_inst : DFF_X1 port map( D => n4247, CK => n828, Q => 
                           REGISTERS_4_63_port, QN => n_1260);
   REGISTERS_reg_4_62_inst : DFF_X1 port map( D => n4246, CK => n828, Q => 
                           REGISTERS_4_62_port, QN => n_1261);
   REGISTERS_reg_4_61_inst : DFF_X1 port map( D => n4245, CK => n828, Q => 
                           REGISTERS_4_61_port, QN => n_1262);
   REGISTERS_reg_4_60_inst : DFF_X1 port map( D => n4244, CK => n828, Q => 
                           REGISTERS_4_60_port, QN => n_1263);
   REGISTERS_reg_4_59_inst : DFF_X1 port map( D => n4243, CK => n828, Q => 
                           REGISTERS_4_59_port, QN => n_1264);
   REGISTERS_reg_4_58_inst : DFF_X1 port map( D => n4242, CK => n828, Q => 
                           REGISTERS_4_58_port, QN => n_1265);
   REGISTERS_reg_4_57_inst : DFF_X1 port map( D => n4241, CK => n828, Q => 
                           REGISTERS_4_57_port, QN => n_1266);
   REGISTERS_reg_4_56_inst : DFF_X1 port map( D => n4240, CK => n828, Q => 
                           REGISTERS_4_56_port, QN => n_1267);
   REGISTERS_reg_4_55_inst : DFF_X1 port map( D => n4239, CK => n828, Q => 
                           REGISTERS_4_55_port, QN => n_1268);
   REGISTERS_reg_4_54_inst : DFF_X1 port map( D => n4238, CK => n828, Q => 
                           REGISTERS_4_54_port, QN => n_1269);
   REGISTERS_reg_4_53_inst : DFF_X1 port map( D => n4237, CK => n828, Q => 
                           REGISTERS_4_53_port, QN => n_1270);
   REGISTERS_reg_4_52_inst : DFF_X1 port map( D => n4236, CK => n829, Q => 
                           REGISTERS_4_52_port, QN => n_1271);
   REGISTERS_reg_4_51_inst : DFF_X1 port map( D => n4235, CK => n829, Q => 
                           REGISTERS_4_51_port, QN => n_1272);
   REGISTERS_reg_4_50_inst : DFF_X1 port map( D => n4234, CK => n829, Q => 
                           REGISTERS_4_50_port, QN => n_1273);
   REGISTERS_reg_4_49_inst : DFF_X1 port map( D => n4233, CK => n829, Q => 
                           REGISTERS_4_49_port, QN => n_1274);
   REGISTERS_reg_4_48_inst : DFF_X1 port map( D => n4232, CK => n829, Q => 
                           REGISTERS_4_48_port, QN => n_1275);
   REGISTERS_reg_4_47_inst : DFF_X1 port map( D => n4231, CK => n829, Q => 
                           REGISTERS_4_47_port, QN => n_1276);
   REGISTERS_reg_4_46_inst : DFF_X1 port map( D => n4230, CK => n829, Q => 
                           REGISTERS_4_46_port, QN => n_1277);
   REGISTERS_reg_4_45_inst : DFF_X1 port map( D => n4229, CK => n829, Q => 
                           REGISTERS_4_45_port, QN => n_1278);
   REGISTERS_reg_4_44_inst : DFF_X1 port map( D => n4228, CK => n829, Q => 
                           REGISTERS_4_44_port, QN => n_1279);
   REGISTERS_reg_4_43_inst : DFF_X1 port map( D => n4227, CK => n829, Q => 
                           REGISTERS_4_43_port, QN => n_1280);
   REGISTERS_reg_4_42_inst : DFF_X1 port map( D => n4226, CK => n829, Q => 
                           REGISTERS_4_42_port, QN => n_1281);
   REGISTERS_reg_4_41_inst : DFF_X1 port map( D => n4225, CK => n830, Q => 
                           REGISTERS_4_41_port, QN => n_1282);
   REGISTERS_reg_4_40_inst : DFF_X1 port map( D => n4224, CK => n830, Q => 
                           REGISTERS_4_40_port, QN => n_1283);
   REGISTERS_reg_4_39_inst : DFF_X1 port map( D => n4223, CK => n830, Q => 
                           REGISTERS_4_39_port, QN => n_1284);
   REGISTERS_reg_4_38_inst : DFF_X1 port map( D => n4222, CK => n830, Q => 
                           REGISTERS_4_38_port, QN => n_1285);
   REGISTERS_reg_4_37_inst : DFF_X1 port map( D => n4221, CK => n830, Q => 
                           REGISTERS_4_37_port, QN => n_1286);
   REGISTERS_reg_4_36_inst : DFF_X1 port map( D => n4220, CK => n830, Q => 
                           REGISTERS_4_36_port, QN => n_1287);
   REGISTERS_reg_4_35_inst : DFF_X1 port map( D => n4219, CK => n830, Q => 
                           REGISTERS_4_35_port, QN => n_1288);
   REGISTERS_reg_4_34_inst : DFF_X1 port map( D => n4218, CK => n830, Q => 
                           REGISTERS_4_34_port, QN => n_1289);
   REGISTERS_reg_4_33_inst : DFF_X1 port map( D => n4217, CK => n830, Q => 
                           REGISTERS_4_33_port, QN => n_1290);
   REGISTERS_reg_4_32_inst : DFF_X1 port map( D => n4216, CK => n830, Q => 
                           REGISTERS_4_32_port, QN => n_1291);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n4215, CK => n830, Q => 
                           REGISTERS_4_31_port, QN => n_1292);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n4214, CK => n831, Q => 
                           REGISTERS_4_30_port, QN => n_1293);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n4213, CK => n831, Q => 
                           REGISTERS_4_29_port, QN => n_1294);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n4212, CK => n831, Q => 
                           REGISTERS_4_28_port, QN => n_1295);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n4211, CK => n831, Q => 
                           REGISTERS_4_27_port, QN => n_1296);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n4210, CK => n831, Q => 
                           REGISTERS_4_26_port, QN => n_1297);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n4209, CK => n831, Q => 
                           REGISTERS_4_25_port, QN => n_1298);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n4208, CK => n831, Q => 
                           REGISTERS_4_24_port, QN => n_1299);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n4207, CK => n831, Q => 
                           REGISTERS_4_23_port, QN => n_1300);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n4206, CK => n831, Q => 
                           REGISTERS_4_22_port, QN => n_1301);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n4205, CK => n831, Q => 
                           REGISTERS_4_21_port, QN => n_1302);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n4204, CK => n831, Q => 
                           REGISTERS_4_20_port, QN => n_1303);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n4203, CK => n832, Q => 
                           REGISTERS_4_19_port, QN => n_1304);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n4202, CK => n832, Q => 
                           REGISTERS_4_18_port, QN => n_1305);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n4201, CK => n832, Q => 
                           REGISTERS_4_17_port, QN => n_1306);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n4200, CK => n832, Q => 
                           REGISTERS_4_16_port, QN => n_1307);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n4199, CK => n832, Q => 
                           REGISTERS_4_15_port, QN => n_1308);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n4198, CK => n832, Q => 
                           REGISTERS_4_14_port, QN => n_1309);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n4197, CK => n832, Q => 
                           REGISTERS_4_13_port, QN => n_1310);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n4196, CK => n832, Q => 
                           REGISTERS_4_12_port, QN => n_1311);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n4195, CK => n832, Q => 
                           REGISTERS_4_11_port, QN => n_1312);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n4194, CK => n832, Q => 
                           REGISTERS_4_10_port, QN => n_1313);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n4193, CK => n832, Q => 
                           REGISTERS_4_9_port, QN => n_1314);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n4192, CK => n833, Q => 
                           REGISTERS_4_8_port, QN => n_1315);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n4191, CK => n833, Q => 
                           REGISTERS_4_7_port, QN => n_1316);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n4190, CK => n833, Q => 
                           REGISTERS_4_6_port, QN => n_1317);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n4189, CK => n833, Q => 
                           REGISTERS_4_5_port, QN => n_1318);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n4188, CK => n833, Q => 
                           REGISTERS_4_4_port, QN => n_1319);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n4187, CK => n833, Q => 
                           REGISTERS_4_3_port, QN => n_1320);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n4186, CK => n833, Q => 
                           REGISTERS_4_2_port, QN => n_1321);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n4185, CK => n833, Q => 
                           REGISTERS_4_1_port, QN => n_1322);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n4184, CK => n833, Q => 
                           REGISTERS_4_0_port, QN => n_1323);
   REGISTERS_reg_5_63_inst : DFF_X1 port map( D => n4183, CK => n833, Q => 
                           REGISTERS_5_63_port, QN => n_1324);
   REGISTERS_reg_5_62_inst : DFF_X1 port map( D => n4182, CK => n833, Q => 
                           REGISTERS_5_62_port, QN => n_1325);
   REGISTERS_reg_5_61_inst : DFF_X1 port map( D => n4181, CK => n834, Q => 
                           REGISTERS_5_61_port, QN => n_1326);
   REGISTERS_reg_5_60_inst : DFF_X1 port map( D => n4180, CK => n834, Q => 
                           REGISTERS_5_60_port, QN => n_1327);
   REGISTERS_reg_5_59_inst : DFF_X1 port map( D => n4179, CK => n834, Q => 
                           REGISTERS_5_59_port, QN => n_1328);
   REGISTERS_reg_5_58_inst : DFF_X1 port map( D => n4178, CK => n834, Q => 
                           REGISTERS_5_58_port, QN => n_1329);
   REGISTERS_reg_5_57_inst : DFF_X1 port map( D => n4177, CK => n834, Q => 
                           REGISTERS_5_57_port, QN => n_1330);
   REGISTERS_reg_5_56_inst : DFF_X1 port map( D => n4176, CK => n834, Q => 
                           REGISTERS_5_56_port, QN => n_1331);
   REGISTERS_reg_5_55_inst : DFF_X1 port map( D => n4175, CK => n834, Q => 
                           REGISTERS_5_55_port, QN => n_1332);
   REGISTERS_reg_5_54_inst : DFF_X1 port map( D => n4174, CK => n834, Q => 
                           REGISTERS_5_54_port, QN => n_1333);
   REGISTERS_reg_5_53_inst : DFF_X1 port map( D => n4173, CK => n834, Q => 
                           REGISTERS_5_53_port, QN => n_1334);
   REGISTERS_reg_5_52_inst : DFF_X1 port map( D => n4172, CK => n834, Q => 
                           REGISTERS_5_52_port, QN => n_1335);
   REGISTERS_reg_5_51_inst : DFF_X1 port map( D => n4171, CK => n834, Q => 
                           REGISTERS_5_51_port, QN => n_1336);
   REGISTERS_reg_5_50_inst : DFF_X1 port map( D => n4170, CK => n835, Q => 
                           REGISTERS_5_50_port, QN => n_1337);
   REGISTERS_reg_5_49_inst : DFF_X1 port map( D => n4169, CK => n835, Q => 
                           REGISTERS_5_49_port, QN => n_1338);
   REGISTERS_reg_5_48_inst : DFF_X1 port map( D => n4168, CK => n835, Q => 
                           REGISTERS_5_48_port, QN => n_1339);
   REGISTERS_reg_5_47_inst : DFF_X1 port map( D => n4167, CK => n835, Q => 
                           REGISTERS_5_47_port, QN => n_1340);
   REGISTERS_reg_5_46_inst : DFF_X1 port map( D => n4166, CK => n835, Q => 
                           REGISTERS_5_46_port, QN => n_1341);
   REGISTERS_reg_5_45_inst : DFF_X1 port map( D => n4165, CK => n835, Q => 
                           REGISTERS_5_45_port, QN => n_1342);
   REGISTERS_reg_5_44_inst : DFF_X1 port map( D => n4164, CK => n835, Q => 
                           REGISTERS_5_44_port, QN => n_1343);
   REGISTERS_reg_5_43_inst : DFF_X1 port map( D => n4163, CK => n835, Q => 
                           REGISTERS_5_43_port, QN => n_1344);
   REGISTERS_reg_5_42_inst : DFF_X1 port map( D => n4162, CK => n835, Q => 
                           REGISTERS_5_42_port, QN => n_1345);
   REGISTERS_reg_5_41_inst : DFF_X1 port map( D => n4161, CK => n835, Q => 
                           REGISTERS_5_41_port, QN => n_1346);
   REGISTERS_reg_5_40_inst : DFF_X1 port map( D => n4160, CK => n835, Q => 
                           REGISTERS_5_40_port, QN => n_1347);
   REGISTERS_reg_5_39_inst : DFF_X1 port map( D => n4159, CK => n836, Q => 
                           REGISTERS_5_39_port, QN => n_1348);
   REGISTERS_reg_5_38_inst : DFF_X1 port map( D => n4158, CK => n836, Q => 
                           REGISTERS_5_38_port, QN => n_1349);
   REGISTERS_reg_5_37_inst : DFF_X1 port map( D => n4157, CK => n836, Q => 
                           REGISTERS_5_37_port, QN => n_1350);
   REGISTERS_reg_5_36_inst : DFF_X1 port map( D => n4156, CK => n836, Q => 
                           REGISTERS_5_36_port, QN => n_1351);
   REGISTERS_reg_5_35_inst : DFF_X1 port map( D => n4155, CK => n836, Q => 
                           REGISTERS_5_35_port, QN => n_1352);
   REGISTERS_reg_5_34_inst : DFF_X1 port map( D => n4154, CK => n836, Q => 
                           REGISTERS_5_34_port, QN => n_1353);
   REGISTERS_reg_5_33_inst : DFF_X1 port map( D => n4153, CK => n836, Q => 
                           REGISTERS_5_33_port, QN => n_1354);
   REGISTERS_reg_5_32_inst : DFF_X1 port map( D => n4152, CK => n836, Q => 
                           REGISTERS_5_32_port, QN => n_1355);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n4151, CK => n836, Q => 
                           REGISTERS_5_31_port, QN => n_1356);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n4150, CK => n836, Q => 
                           REGISTERS_5_30_port, QN => n_1357);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n4149, CK => n836, Q => 
                           REGISTERS_5_29_port, QN => n_1358);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n4148, CK => n837, Q => 
                           REGISTERS_5_28_port, QN => n_1359);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n4147, CK => n837, Q => 
                           REGISTERS_5_27_port, QN => n_1360);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n4146, CK => n837, Q => 
                           REGISTERS_5_26_port, QN => n_1361);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n4145, CK => n837, Q => 
                           REGISTERS_5_25_port, QN => n_1362);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n4144, CK => n837, Q => 
                           REGISTERS_5_24_port, QN => n_1363);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n4143, CK => n837, Q => 
                           REGISTERS_5_23_port, QN => n_1364);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n4142, CK => n837, Q => 
                           REGISTERS_5_22_port, QN => n_1365);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n4141, CK => n837, Q => 
                           REGISTERS_5_21_port, QN => n_1366);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n4140, CK => n837, Q => 
                           REGISTERS_5_20_port, QN => n_1367);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n4139, CK => n837, Q => 
                           REGISTERS_5_19_port, QN => n_1368);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n4138, CK => n837, Q => 
                           REGISTERS_5_18_port, QN => n_1369);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n4137, CK => n838, Q => 
                           REGISTERS_5_17_port, QN => n_1370);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n4136, CK => n838, Q => 
                           REGISTERS_5_16_port, QN => n_1371);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n4135, CK => n838, Q => 
                           REGISTERS_5_15_port, QN => n_1372);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n4134, CK => n838, Q => 
                           REGISTERS_5_14_port, QN => n_1373);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n4133, CK => n838, Q => 
                           REGISTERS_5_13_port, QN => n_1374);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n4132, CK => n838, Q => 
                           REGISTERS_5_12_port, QN => n_1375);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n4131, CK => n838, Q => 
                           REGISTERS_5_11_port, QN => n_1376);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n4130, CK => n838, Q => 
                           REGISTERS_5_10_port, QN => n_1377);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n4129, CK => n838, Q => 
                           REGISTERS_5_9_port, QN => n_1378);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n4128, CK => n838, Q => 
                           REGISTERS_5_8_port, QN => n_1379);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n4127, CK => n838, Q => 
                           REGISTERS_5_7_port, QN => n_1380);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n4126, CK => n839, Q => 
                           REGISTERS_5_6_port, QN => n_1381);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n4125, CK => n839, Q => 
                           REGISTERS_5_5_port, QN => n_1382);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n4124, CK => n839, Q => 
                           REGISTERS_5_4_port, QN => n_1383);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n4123, CK => n839, Q => 
                           REGISTERS_5_3_port, QN => n_1384);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n4122, CK => n839, Q => 
                           REGISTERS_5_2_port, QN => n_1385);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n4121, CK => n839, Q => 
                           REGISTERS_5_1_port, QN => n_1386);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n4120, CK => n839, Q => 
                           REGISTERS_5_0_port, QN => n_1387);
   REGISTERS_reg_6_63_inst : DFF_X1 port map( D => n4119, CK => n839, Q => 
                           REGISTERS_6_63_port, QN => n_1388);
   REGISTERS_reg_6_62_inst : DFF_X1 port map( D => n4118, CK => n839, Q => 
                           REGISTERS_6_62_port, QN => n_1389);
   REGISTERS_reg_6_61_inst : DFF_X1 port map( D => n4117, CK => n839, Q => 
                           REGISTERS_6_61_port, QN => n_1390);
   REGISTERS_reg_6_60_inst : DFF_X1 port map( D => n4116, CK => n839, Q => 
                           REGISTERS_6_60_port, QN => n_1391);
   REGISTERS_reg_6_59_inst : DFF_X1 port map( D => n4115, CK => n840, Q => 
                           REGISTERS_6_59_port, QN => n_1392);
   REGISTERS_reg_6_58_inst : DFF_X1 port map( D => n4114, CK => n840, Q => 
                           REGISTERS_6_58_port, QN => n_1393);
   REGISTERS_reg_6_57_inst : DFF_X1 port map( D => n4113, CK => n840, Q => 
                           REGISTERS_6_57_port, QN => n_1394);
   REGISTERS_reg_6_56_inst : DFF_X1 port map( D => n4112, CK => n840, Q => 
                           REGISTERS_6_56_port, QN => n_1395);
   REGISTERS_reg_6_55_inst : DFF_X1 port map( D => n4111, CK => n840, Q => 
                           REGISTERS_6_55_port, QN => n_1396);
   REGISTERS_reg_6_54_inst : DFF_X1 port map( D => n4110, CK => n840, Q => 
                           REGISTERS_6_54_port, QN => n_1397);
   REGISTERS_reg_6_53_inst : DFF_X1 port map( D => n4109, CK => n840, Q => 
                           REGISTERS_6_53_port, QN => n_1398);
   REGISTERS_reg_6_52_inst : DFF_X1 port map( D => n4108, CK => n840, Q => 
                           REGISTERS_6_52_port, QN => n_1399);
   REGISTERS_reg_6_51_inst : DFF_X1 port map( D => n4107, CK => n840, Q => 
                           REGISTERS_6_51_port, QN => n_1400);
   REGISTERS_reg_6_50_inst : DFF_X1 port map( D => n4106, CK => n840, Q => 
                           REGISTERS_6_50_port, QN => n_1401);
   REGISTERS_reg_6_49_inst : DFF_X1 port map( D => n4105, CK => n840, Q => 
                           REGISTERS_6_49_port, QN => n_1402);
   REGISTERS_reg_6_48_inst : DFF_X1 port map( D => n4104, CK => n841, Q => 
                           REGISTERS_6_48_port, QN => n_1403);
   REGISTERS_reg_6_47_inst : DFF_X1 port map( D => n4103, CK => n841, Q => 
                           REGISTERS_6_47_port, QN => n_1404);
   REGISTERS_reg_6_46_inst : DFF_X1 port map( D => n4102, CK => n841, Q => 
                           REGISTERS_6_46_port, QN => n_1405);
   REGISTERS_reg_6_45_inst : DFF_X1 port map( D => n4101, CK => n841, Q => 
                           REGISTERS_6_45_port, QN => n_1406);
   REGISTERS_reg_6_44_inst : DFF_X1 port map( D => n4100, CK => n841, Q => 
                           REGISTERS_6_44_port, QN => n_1407);
   REGISTERS_reg_6_43_inst : DFF_X1 port map( D => n4099, CK => n841, Q => 
                           REGISTERS_6_43_port, QN => n_1408);
   REGISTERS_reg_6_42_inst : DFF_X1 port map( D => n4098, CK => n841, Q => 
                           REGISTERS_6_42_port, QN => n_1409);
   REGISTERS_reg_6_41_inst : DFF_X1 port map( D => n4097, CK => n841, Q => 
                           REGISTERS_6_41_port, QN => n_1410);
   REGISTERS_reg_6_40_inst : DFF_X1 port map( D => n4096, CK => n841, Q => 
                           REGISTERS_6_40_port, QN => n_1411);
   REGISTERS_reg_6_39_inst : DFF_X1 port map( D => n4095, CK => n841, Q => 
                           REGISTERS_6_39_port, QN => n_1412);
   REGISTERS_reg_6_38_inst : DFF_X1 port map( D => n4094, CK => n841, Q => 
                           REGISTERS_6_38_port, QN => n_1413);
   REGISTERS_reg_6_37_inst : DFF_X1 port map( D => n4093, CK => n842, Q => 
                           REGISTERS_6_37_port, QN => n_1414);
   REGISTERS_reg_6_36_inst : DFF_X1 port map( D => n4092, CK => n842, Q => 
                           REGISTERS_6_36_port, QN => n_1415);
   REGISTERS_reg_6_35_inst : DFF_X1 port map( D => n4091, CK => n842, Q => 
                           REGISTERS_6_35_port, QN => n_1416);
   REGISTERS_reg_6_34_inst : DFF_X1 port map( D => n4090, CK => n842, Q => 
                           REGISTERS_6_34_port, QN => n_1417);
   REGISTERS_reg_6_33_inst : DFF_X1 port map( D => n4089, CK => n842, Q => 
                           REGISTERS_6_33_port, QN => n_1418);
   REGISTERS_reg_6_32_inst : DFF_X1 port map( D => n4088, CK => n842, Q => 
                           REGISTERS_6_32_port, QN => n_1419);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n4087, CK => n842, Q => 
                           REGISTERS_6_31_port, QN => n_1420);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n4086, CK => n842, Q => 
                           REGISTERS_6_30_port, QN => n_1421);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n4085, CK => n842, Q => 
                           REGISTERS_6_29_port, QN => n_1422);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n4084, CK => n842, Q => 
                           REGISTERS_6_28_port, QN => n_1423);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n4083, CK => n842, Q => 
                           REGISTERS_6_27_port, QN => n_1424);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n4082, CK => n843, Q => 
                           REGISTERS_6_26_port, QN => n_1425);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n4081, CK => n843, Q => 
                           REGISTERS_6_25_port, QN => n_1426);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n4080, CK => n843, Q => 
                           REGISTERS_6_24_port, QN => n_1427);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n4079, CK => n843, Q => 
                           REGISTERS_6_23_port, QN => n_1428);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n4078, CK => n843, Q => 
                           REGISTERS_6_22_port, QN => n_1429);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n4077, CK => n843, Q => 
                           REGISTERS_6_21_port, QN => n_1430);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n4076, CK => n843, Q => 
                           REGISTERS_6_20_port, QN => n_1431);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n4075, CK => n843, Q => 
                           REGISTERS_6_19_port, QN => n_1432);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n4074, CK => n843, Q => 
                           REGISTERS_6_18_port, QN => n_1433);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n4073, CK => n843, Q => 
                           REGISTERS_6_17_port, QN => n_1434);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n4072, CK => n843, Q => 
                           REGISTERS_6_16_port, QN => n_1435);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n4071, CK => n844, Q => 
                           REGISTERS_6_15_port, QN => n_1436);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n4070, CK => n844, Q => 
                           REGISTERS_6_14_port, QN => n_1437);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n4069, CK => n844, Q => 
                           REGISTERS_6_13_port, QN => n_1438);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n4068, CK => n844, Q => 
                           REGISTERS_6_12_port, QN => n_1439);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n4067, CK => n844, Q => 
                           REGISTERS_6_11_port, QN => n_1440);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n4066, CK => n844, Q => 
                           REGISTERS_6_10_port, QN => n_1441);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n4065, CK => n844, Q => 
                           REGISTERS_6_9_port, QN => n_1442);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n4064, CK => n844, Q => 
                           REGISTERS_6_8_port, QN => n_1443);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n4063, CK => n844, Q => 
                           REGISTERS_6_7_port, QN => n_1444);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n4062, CK => n844, Q => 
                           REGISTERS_6_6_port, QN => n_1445);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n4061, CK => n844, Q => 
                           REGISTERS_6_5_port, QN => n_1446);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n4060, CK => n845, Q => 
                           REGISTERS_6_4_port, QN => n_1447);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n4059, CK => n845, Q => 
                           REGISTERS_6_3_port, QN => n_1448);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n4058, CK => n845, Q => 
                           REGISTERS_6_2_port, QN => n_1449);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n4057, CK => n845, Q => 
                           REGISTERS_6_1_port, QN => n_1450);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n4056, CK => n845, Q => 
                           REGISTERS_6_0_port, QN => n_1451);
   REGISTERS_reg_7_63_inst : DFF_X1 port map( D => n4055, CK => n845, Q => 
                           REGISTERS_7_63_port, QN => n_1452);
   REGISTERS_reg_7_62_inst : DFF_X1 port map( D => n4054, CK => n845, Q => 
                           REGISTERS_7_62_port, QN => n_1453);
   REGISTERS_reg_7_61_inst : DFF_X1 port map( D => n4053, CK => n845, Q => 
                           REGISTERS_7_61_port, QN => n_1454);
   REGISTERS_reg_7_60_inst : DFF_X1 port map( D => n4052, CK => n845, Q => 
                           REGISTERS_7_60_port, QN => n_1455);
   REGISTERS_reg_7_59_inst : DFF_X1 port map( D => n4051, CK => n845, Q => 
                           REGISTERS_7_59_port, QN => n_1456);
   REGISTERS_reg_7_58_inst : DFF_X1 port map( D => n4050, CK => n845, Q => 
                           REGISTERS_7_58_port, QN => n_1457);
   REGISTERS_reg_7_57_inst : DFF_X1 port map( D => n4049, CK => n846, Q => 
                           REGISTERS_7_57_port, QN => n_1458);
   REGISTERS_reg_7_56_inst : DFF_X1 port map( D => n4048, CK => n846, Q => 
                           REGISTERS_7_56_port, QN => n_1459);
   REGISTERS_reg_7_55_inst : DFF_X1 port map( D => n4047, CK => n846, Q => 
                           REGISTERS_7_55_port, QN => n_1460);
   REGISTERS_reg_7_54_inst : DFF_X1 port map( D => n4046, CK => n846, Q => 
                           REGISTERS_7_54_port, QN => n_1461);
   REGISTERS_reg_7_53_inst : DFF_X1 port map( D => n4045, CK => n846, Q => 
                           REGISTERS_7_53_port, QN => n_1462);
   REGISTERS_reg_7_52_inst : DFF_X1 port map( D => n4044, CK => n846, Q => 
                           REGISTERS_7_52_port, QN => n_1463);
   REGISTERS_reg_7_51_inst : DFF_X1 port map( D => n4043, CK => n846, Q => 
                           REGISTERS_7_51_port, QN => n_1464);
   REGISTERS_reg_7_50_inst : DFF_X1 port map( D => n4042, CK => n846, Q => 
                           REGISTERS_7_50_port, QN => n_1465);
   REGISTERS_reg_7_49_inst : DFF_X1 port map( D => n4041, CK => n846, Q => 
                           REGISTERS_7_49_port, QN => n_1466);
   REGISTERS_reg_7_48_inst : DFF_X1 port map( D => n4040, CK => n846, Q => 
                           REGISTERS_7_48_port, QN => n_1467);
   REGISTERS_reg_7_47_inst : DFF_X1 port map( D => n4039, CK => n846, Q => 
                           REGISTERS_7_47_port, QN => n_1468);
   REGISTERS_reg_7_46_inst : DFF_X1 port map( D => n4038, CK => n847, Q => 
                           REGISTERS_7_46_port, QN => n_1469);
   REGISTERS_reg_7_45_inst : DFF_X1 port map( D => n4037, CK => n847, Q => 
                           REGISTERS_7_45_port, QN => n_1470);
   REGISTERS_reg_7_44_inst : DFF_X1 port map( D => n4036, CK => n847, Q => 
                           REGISTERS_7_44_port, QN => n_1471);
   REGISTERS_reg_7_43_inst : DFF_X1 port map( D => n4035, CK => n847, Q => 
                           REGISTERS_7_43_port, QN => n_1472);
   REGISTERS_reg_7_42_inst : DFF_X1 port map( D => n4034, CK => n847, Q => 
                           REGISTERS_7_42_port, QN => n_1473);
   REGISTERS_reg_7_41_inst : DFF_X1 port map( D => n4033, CK => n847, Q => 
                           REGISTERS_7_41_port, QN => n_1474);
   REGISTERS_reg_7_40_inst : DFF_X1 port map( D => n4032, CK => n847, Q => 
                           REGISTERS_7_40_port, QN => n_1475);
   REGISTERS_reg_7_39_inst : DFF_X1 port map( D => n4031, CK => n847, Q => 
                           REGISTERS_7_39_port, QN => n_1476);
   REGISTERS_reg_7_38_inst : DFF_X1 port map( D => n4030, CK => n847, Q => 
                           REGISTERS_7_38_port, QN => n_1477);
   REGISTERS_reg_7_37_inst : DFF_X1 port map( D => n4029, CK => n847, Q => 
                           REGISTERS_7_37_port, QN => n_1478);
   REGISTERS_reg_7_36_inst : DFF_X1 port map( D => n4028, CK => n847, Q => 
                           REGISTERS_7_36_port, QN => n_1479);
   REGISTERS_reg_7_35_inst : DFF_X1 port map( D => n4027, CK => n848, Q => 
                           REGISTERS_7_35_port, QN => n_1480);
   REGISTERS_reg_7_34_inst : DFF_X1 port map( D => n4026, CK => n848, Q => 
                           REGISTERS_7_34_port, QN => n_1481);
   REGISTERS_reg_7_33_inst : DFF_X1 port map( D => n4025, CK => n848, Q => 
                           REGISTERS_7_33_port, QN => n_1482);
   REGISTERS_reg_7_32_inst : DFF_X1 port map( D => n4024, CK => n848, Q => 
                           REGISTERS_7_32_port, QN => n_1483);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n4023, CK => n848, Q => 
                           REGISTERS_7_31_port, QN => n_1484);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n4022, CK => n848, Q => 
                           REGISTERS_7_30_port, QN => n_1485);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n4021, CK => n848, Q => 
                           REGISTERS_7_29_port, QN => n_1486);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n4020, CK => n848, Q => 
                           REGISTERS_7_28_port, QN => n_1487);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n4019, CK => n848, Q => 
                           REGISTERS_7_27_port, QN => n_1488);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n4018, CK => n848, Q => 
                           REGISTERS_7_26_port, QN => n_1489);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n4017, CK => n848, Q => 
                           REGISTERS_7_25_port, QN => n_1490);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n4016, CK => n849, Q => 
                           REGISTERS_7_24_port, QN => n_1491);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n4015, CK => n849, Q => 
                           REGISTERS_7_23_port, QN => n_1492);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n4014, CK => n849, Q => 
                           REGISTERS_7_22_port, QN => n_1493);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n4013, CK => n849, Q => 
                           REGISTERS_7_21_port, QN => n_1494);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n4012, CK => n849, Q => 
                           REGISTERS_7_20_port, QN => n_1495);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n4011, CK => n849, Q => 
                           REGISTERS_7_19_port, QN => n_1496);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n4010, CK => n849, Q => 
                           REGISTERS_7_18_port, QN => n_1497);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n4009, CK => n849, Q => 
                           REGISTERS_7_17_port, QN => n_1498);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n4008, CK => n849, Q => 
                           REGISTERS_7_16_port, QN => n_1499);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n4007, CK => n849, Q => 
                           REGISTERS_7_15_port, QN => n_1500);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n4006, CK => n849, Q => 
                           REGISTERS_7_14_port, QN => n_1501);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n4005, CK => n850, Q => 
                           REGISTERS_7_13_port, QN => n_1502);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n4004, CK => n850, Q => 
                           REGISTERS_7_12_port, QN => n_1503);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n4003, CK => n850, Q => 
                           REGISTERS_7_11_port, QN => n_1504);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n4002, CK => n850, Q => 
                           REGISTERS_7_10_port, QN => n_1505);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n4001, CK => n850, Q => 
                           REGISTERS_7_9_port, QN => n_1506);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n4000, CK => n850, Q => 
                           REGISTERS_7_8_port, QN => n_1507);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n3999, CK => n850, Q => 
                           REGISTERS_7_7_port, QN => n_1508);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n3998, CK => n850, Q => 
                           REGISTERS_7_6_port, QN => n_1509);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n3997, CK => n850, Q => 
                           REGISTERS_7_5_port, QN => n_1510);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n3996, CK => n850, Q => 
                           REGISTERS_7_4_port, QN => n_1511);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n3995, CK => n850, Q => 
                           REGISTERS_7_3_port, QN => n_1512);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n3994, CK => n851, Q => 
                           REGISTERS_7_2_port, QN => n_1513);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n3993, CK => n851, Q => 
                           REGISTERS_7_1_port, QN => n_1514);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n3992, CK => n851, Q => 
                           REGISTERS_7_0_port, QN => n_1515);
   REGISTERS_reg_8_63_inst : DFF_X1 port map( D => n3991, CK => n851, Q => 
                           REGISTERS_8_63_port, QN => n_1516);
   REGISTERS_reg_8_62_inst : DFF_X1 port map( D => n3990, CK => n851, Q => 
                           REGISTERS_8_62_port, QN => n_1517);
   REGISTERS_reg_8_61_inst : DFF_X1 port map( D => n3989, CK => n851, Q => 
                           REGISTERS_8_61_port, QN => n_1518);
   REGISTERS_reg_8_60_inst : DFF_X1 port map( D => n3988, CK => n851, Q => 
                           REGISTERS_8_60_port, QN => n_1519);
   REGISTERS_reg_8_59_inst : DFF_X1 port map( D => n3987, CK => n851, Q => 
                           REGISTERS_8_59_port, QN => n_1520);
   REGISTERS_reg_8_58_inst : DFF_X1 port map( D => n3986, CK => n851, Q => 
                           REGISTERS_8_58_port, QN => n_1521);
   REGISTERS_reg_8_57_inst : DFF_X1 port map( D => n3985, CK => n851, Q => 
                           REGISTERS_8_57_port, QN => n_1522);
   REGISTERS_reg_8_56_inst : DFF_X1 port map( D => n3984, CK => n851, Q => 
                           REGISTERS_8_56_port, QN => n_1523);
   REGISTERS_reg_8_55_inst : DFF_X1 port map( D => n3983, CK => n852, Q => 
                           REGISTERS_8_55_port, QN => n_1524);
   REGISTERS_reg_8_54_inst : DFF_X1 port map( D => n3982, CK => n852, Q => 
                           REGISTERS_8_54_port, QN => n_1525);
   REGISTERS_reg_8_53_inst : DFF_X1 port map( D => n3981, CK => n852, Q => 
                           REGISTERS_8_53_port, QN => n_1526);
   REGISTERS_reg_8_52_inst : DFF_X1 port map( D => n3980, CK => n852, Q => 
                           REGISTERS_8_52_port, QN => n_1527);
   REGISTERS_reg_8_51_inst : DFF_X1 port map( D => n3979, CK => n852, Q => 
                           REGISTERS_8_51_port, QN => n_1528);
   REGISTERS_reg_8_50_inst : DFF_X1 port map( D => n3978, CK => n852, Q => 
                           REGISTERS_8_50_port, QN => n_1529);
   REGISTERS_reg_8_49_inst : DFF_X1 port map( D => n3977, CK => n852, Q => 
                           REGISTERS_8_49_port, QN => n_1530);
   REGISTERS_reg_8_48_inst : DFF_X1 port map( D => n3976, CK => n852, Q => 
                           REGISTERS_8_48_port, QN => n_1531);
   REGISTERS_reg_8_47_inst : DFF_X1 port map( D => n3975, CK => n852, Q => 
                           REGISTERS_8_47_port, QN => n_1532);
   REGISTERS_reg_8_46_inst : DFF_X1 port map( D => n3974, CK => n852, Q => 
                           REGISTERS_8_46_port, QN => n_1533);
   REGISTERS_reg_8_45_inst : DFF_X1 port map( D => n3973, CK => n852, Q => 
                           REGISTERS_8_45_port, QN => n_1534);
   REGISTERS_reg_8_44_inst : DFF_X1 port map( D => n3972, CK => n853, Q => 
                           REGISTERS_8_44_port, QN => n_1535);
   REGISTERS_reg_8_43_inst : DFF_X1 port map( D => n3971, CK => n853, Q => 
                           REGISTERS_8_43_port, QN => n_1536);
   REGISTERS_reg_8_42_inst : DFF_X1 port map( D => n3970, CK => n853, Q => 
                           REGISTERS_8_42_port, QN => n_1537);
   REGISTERS_reg_8_41_inst : DFF_X1 port map( D => n3969, CK => n853, Q => 
                           REGISTERS_8_41_port, QN => n_1538);
   REGISTERS_reg_8_40_inst : DFF_X1 port map( D => n3968, CK => n853, Q => 
                           REGISTERS_8_40_port, QN => n_1539);
   REGISTERS_reg_8_39_inst : DFF_X1 port map( D => n3967, CK => n853, Q => 
                           REGISTERS_8_39_port, QN => n_1540);
   REGISTERS_reg_8_38_inst : DFF_X1 port map( D => n3966, CK => n853, Q => 
                           REGISTERS_8_38_port, QN => n_1541);
   REGISTERS_reg_8_37_inst : DFF_X1 port map( D => n3965, CK => n853, Q => 
                           REGISTERS_8_37_port, QN => n_1542);
   REGISTERS_reg_8_36_inst : DFF_X1 port map( D => n3964, CK => n853, Q => 
                           REGISTERS_8_36_port, QN => n_1543);
   REGISTERS_reg_8_35_inst : DFF_X1 port map( D => n3963, CK => n853, Q => 
                           REGISTERS_8_35_port, QN => n_1544);
   REGISTERS_reg_8_34_inst : DFF_X1 port map( D => n3962, CK => n853, Q => 
                           REGISTERS_8_34_port, QN => n_1545);
   REGISTERS_reg_8_33_inst : DFF_X1 port map( D => n3961, CK => n854, Q => 
                           REGISTERS_8_33_port, QN => n_1546);
   REGISTERS_reg_8_32_inst : DFF_X1 port map( D => n3960, CK => n854, Q => 
                           REGISTERS_8_32_port, QN => n_1547);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n3959, CK => n854, Q => 
                           REGISTERS_8_31_port, QN => n_1548);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n3958, CK => n854, Q => 
                           REGISTERS_8_30_port, QN => n_1549);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n3957, CK => n854, Q => 
                           REGISTERS_8_29_port, QN => n_1550);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n3956, CK => n854, Q => 
                           REGISTERS_8_28_port, QN => n_1551);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n3955, CK => n854, Q => 
                           REGISTERS_8_27_port, QN => n_1552);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n3954, CK => n854, Q => 
                           REGISTERS_8_26_port, QN => n_1553);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n3953, CK => n854, Q => 
                           REGISTERS_8_25_port, QN => n_1554);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n3952, CK => n854, Q => 
                           REGISTERS_8_24_port, QN => n_1555);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n3951, CK => n854, Q => 
                           REGISTERS_8_23_port, QN => n_1556);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n3950, CK => n855, Q => 
                           REGISTERS_8_22_port, QN => n_1557);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n3949, CK => n855, Q => 
                           REGISTERS_8_21_port, QN => n_1558);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n3948, CK => n855, Q => 
                           REGISTERS_8_20_port, QN => n_1559);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n3947, CK => n855, Q => 
                           REGISTERS_8_19_port, QN => n_1560);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n3946, CK => n855, Q => 
                           REGISTERS_8_18_port, QN => n_1561);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n3945, CK => n855, Q => 
                           REGISTERS_8_17_port, QN => n_1562);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n3944, CK => n855, Q => 
                           REGISTERS_8_16_port, QN => n_1563);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n3943, CK => n855, Q => 
                           REGISTERS_8_15_port, QN => n_1564);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n3942, CK => n855, Q => 
                           REGISTERS_8_14_port, QN => n_1565);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n3941, CK => n855, Q => 
                           REGISTERS_8_13_port, QN => n_1566);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n3940, CK => n855, Q => 
                           REGISTERS_8_12_port, QN => n_1567);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n3939, CK => n856, Q => 
                           REGISTERS_8_11_port, QN => n_1568);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n3938, CK => n856, Q => 
                           REGISTERS_8_10_port, QN => n_1569);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n3937, CK => n856, Q => 
                           REGISTERS_8_9_port, QN => n_1570);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n3936, CK => n856, Q => 
                           REGISTERS_8_8_port, QN => n_1571);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n3935, CK => n856, Q => 
                           REGISTERS_8_7_port, QN => n_1572);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n3934, CK => n856, Q => 
                           REGISTERS_8_6_port, QN => n_1573);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n3933, CK => n856, Q => 
                           REGISTERS_8_5_port, QN => n_1574);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n3932, CK => n856, Q => 
                           REGISTERS_8_4_port, QN => n_1575);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n3931, CK => n856, Q => 
                           REGISTERS_8_3_port, QN => n_1576);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n3930, CK => n856, Q => 
                           REGISTERS_8_2_port, QN => n_1577);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n3929, CK => n856, Q => 
                           REGISTERS_8_1_port, QN => n_1578);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n3928, CK => n857, Q => 
                           REGISTERS_8_0_port, QN => n_1579);
   REGISTERS_reg_9_63_inst : DFF_X1 port map( D => n3927, CK => n857, Q => 
                           REGISTERS_9_63_port, QN => n_1580);
   REGISTERS_reg_9_62_inst : DFF_X1 port map( D => n3926, CK => n857, Q => 
                           REGISTERS_9_62_port, QN => n_1581);
   REGISTERS_reg_9_61_inst : DFF_X1 port map( D => n3925, CK => n857, Q => 
                           REGISTERS_9_61_port, QN => n_1582);
   REGISTERS_reg_9_60_inst : DFF_X1 port map( D => n3924, CK => n857, Q => 
                           REGISTERS_9_60_port, QN => n_1583);
   REGISTERS_reg_9_59_inst : DFF_X1 port map( D => n3923, CK => n857, Q => 
                           REGISTERS_9_59_port, QN => n_1584);
   REGISTERS_reg_9_58_inst : DFF_X1 port map( D => n3922, CK => n857, Q => 
                           REGISTERS_9_58_port, QN => n_1585);
   REGISTERS_reg_9_57_inst : DFF_X1 port map( D => n3921, CK => n857, Q => 
                           REGISTERS_9_57_port, QN => n_1586);
   REGISTERS_reg_9_56_inst : DFF_X1 port map( D => n3920, CK => n857, Q => 
                           REGISTERS_9_56_port, QN => n_1587);
   REGISTERS_reg_9_55_inst : DFF_X1 port map( D => n3919, CK => n857, Q => 
                           REGISTERS_9_55_port, QN => n_1588);
   REGISTERS_reg_9_54_inst : DFF_X1 port map( D => n3918, CK => n857, Q => 
                           REGISTERS_9_54_port, QN => n_1589);
   REGISTERS_reg_9_53_inst : DFF_X1 port map( D => n3917, CK => n858, Q => 
                           REGISTERS_9_53_port, QN => n_1590);
   REGISTERS_reg_9_52_inst : DFF_X1 port map( D => n3916, CK => n858, Q => 
                           REGISTERS_9_52_port, QN => n_1591);
   REGISTERS_reg_9_51_inst : DFF_X1 port map( D => n3915, CK => n858, Q => 
                           REGISTERS_9_51_port, QN => n_1592);
   REGISTERS_reg_9_50_inst : DFF_X1 port map( D => n3914, CK => n858, Q => 
                           REGISTERS_9_50_port, QN => n_1593);
   REGISTERS_reg_9_49_inst : DFF_X1 port map( D => n3913, CK => n858, Q => 
                           REGISTERS_9_49_port, QN => n_1594);
   REGISTERS_reg_9_48_inst : DFF_X1 port map( D => n3912, CK => n858, Q => 
                           REGISTERS_9_48_port, QN => n_1595);
   REGISTERS_reg_9_47_inst : DFF_X1 port map( D => n3911, CK => n858, Q => 
                           REGISTERS_9_47_port, QN => n_1596);
   REGISTERS_reg_9_46_inst : DFF_X1 port map( D => n3910, CK => n858, Q => 
                           REGISTERS_9_46_port, QN => n_1597);
   REGISTERS_reg_9_45_inst : DFF_X1 port map( D => n3909, CK => n858, Q => 
                           REGISTERS_9_45_port, QN => n_1598);
   REGISTERS_reg_9_44_inst : DFF_X1 port map( D => n3908, CK => n858, Q => 
                           REGISTERS_9_44_port, QN => n_1599);
   REGISTERS_reg_9_43_inst : DFF_X1 port map( D => n3907, CK => n858, Q => 
                           REGISTERS_9_43_port, QN => n_1600);
   REGISTERS_reg_9_42_inst : DFF_X1 port map( D => n3906, CK => n859, Q => 
                           REGISTERS_9_42_port, QN => n_1601);
   REGISTERS_reg_9_41_inst : DFF_X1 port map( D => n3905, CK => n859, Q => 
                           REGISTERS_9_41_port, QN => n_1602);
   REGISTERS_reg_9_40_inst : DFF_X1 port map( D => n3904, CK => n859, Q => 
                           REGISTERS_9_40_port, QN => n_1603);
   REGISTERS_reg_9_39_inst : DFF_X1 port map( D => n3903, CK => n859, Q => 
                           REGISTERS_9_39_port, QN => n_1604);
   REGISTERS_reg_9_38_inst : DFF_X1 port map( D => n3902, CK => n859, Q => 
                           REGISTERS_9_38_port, QN => n_1605);
   REGISTERS_reg_9_37_inst : DFF_X1 port map( D => n3901, CK => n859, Q => 
                           REGISTERS_9_37_port, QN => n_1606);
   REGISTERS_reg_9_36_inst : DFF_X1 port map( D => n3900, CK => n859, Q => 
                           REGISTERS_9_36_port, QN => n_1607);
   REGISTERS_reg_9_35_inst : DFF_X1 port map( D => n3899, CK => n859, Q => 
                           REGISTERS_9_35_port, QN => n_1608);
   REGISTERS_reg_9_34_inst : DFF_X1 port map( D => n3898, CK => n859, Q => 
                           REGISTERS_9_34_port, QN => n_1609);
   REGISTERS_reg_9_33_inst : DFF_X1 port map( D => n3897, CK => n859, Q => 
                           REGISTERS_9_33_port, QN => n_1610);
   REGISTERS_reg_9_32_inst : DFF_X1 port map( D => n3896, CK => n859, Q => 
                           REGISTERS_9_32_port, QN => n_1611);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n3895, CK => n860, Q => 
                           REGISTERS_9_31_port, QN => n_1612);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n3894, CK => n860, Q => 
                           REGISTERS_9_30_port, QN => n_1613);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n3893, CK => n860, Q => 
                           REGISTERS_9_29_port, QN => n_1614);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n3892, CK => n860, Q => 
                           REGISTERS_9_28_port, QN => n_1615);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n3891, CK => n860, Q => 
                           REGISTERS_9_27_port, QN => n_1616);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n3890, CK => n860, Q => 
                           REGISTERS_9_26_port, QN => n_1617);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n3889, CK => n860, Q => 
                           REGISTERS_9_25_port, QN => n_1618);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n3888, CK => n860, Q => 
                           REGISTERS_9_24_port, QN => n_1619);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n3887, CK => n860, Q => 
                           REGISTERS_9_23_port, QN => n_1620);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n3886, CK => n860, Q => 
                           REGISTERS_9_22_port, QN => n_1621);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n3885, CK => n860, Q => 
                           REGISTERS_9_21_port, QN => n_1622);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n3884, CK => n861, Q => 
                           REGISTERS_9_20_port, QN => n_1623);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n3883, CK => n861, Q => 
                           REGISTERS_9_19_port, QN => n_1624);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n3882, CK => n861, Q => 
                           REGISTERS_9_18_port, QN => n_1625);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n3881, CK => n861, Q => 
                           REGISTERS_9_17_port, QN => n_1626);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n3880, CK => n861, Q => 
                           REGISTERS_9_16_port, QN => n_1627);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n3879, CK => n861, Q => 
                           REGISTERS_9_15_port, QN => n_1628);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n3878, CK => n861, Q => 
                           REGISTERS_9_14_port, QN => n_1629);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n3877, CK => n861, Q => 
                           REGISTERS_9_13_port, QN => n_1630);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n3876, CK => n861, Q => 
                           REGISTERS_9_12_port, QN => n_1631);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n3875, CK => n861, Q => 
                           REGISTERS_9_11_port, QN => n_1632);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n3874, CK => n861, Q => 
                           REGISTERS_9_10_port, QN => n_1633);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n3873, CK => n862, Q => 
                           REGISTERS_9_9_port, QN => n_1634);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n3872, CK => n862, Q => 
                           REGISTERS_9_8_port, QN => n_1635);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n3871, CK => n862, Q => 
                           REGISTERS_9_7_port, QN => n_1636);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n3870, CK => n862, Q => 
                           REGISTERS_9_6_port, QN => n_1637);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n3869, CK => n862, Q => 
                           REGISTERS_9_5_port, QN => n_1638);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n3868, CK => n862, Q => 
                           REGISTERS_9_4_port, QN => n_1639);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n3867, CK => n862, Q => 
                           REGISTERS_9_3_port, QN => n_1640);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n3866, CK => n862, Q => 
                           REGISTERS_9_2_port, QN => n_1641);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n3865, CK => n862, Q => 
                           REGISTERS_9_1_port, QN => n_1642);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n3864, CK => n862, Q => 
                           REGISTERS_9_0_port, QN => n_1643);
   REGISTERS_reg_10_63_inst : DFF_X1 port map( D => n3863, CK => n862, Q => 
                           REGISTERS_10_63_port, QN => n_1644);
   REGISTERS_reg_10_62_inst : DFF_X1 port map( D => n3862, CK => n863, Q => 
                           REGISTERS_10_62_port, QN => n_1645);
   REGISTERS_reg_10_61_inst : DFF_X1 port map( D => n3861, CK => n863, Q => 
                           REGISTERS_10_61_port, QN => n_1646);
   REGISTERS_reg_10_60_inst : DFF_X1 port map( D => n3860, CK => n863, Q => 
                           REGISTERS_10_60_port, QN => n_1647);
   REGISTERS_reg_10_59_inst : DFF_X1 port map( D => n3859, CK => n863, Q => 
                           REGISTERS_10_59_port, QN => n_1648);
   REGISTERS_reg_10_58_inst : DFF_X1 port map( D => n3858, CK => n863, Q => 
                           REGISTERS_10_58_port, QN => n_1649);
   REGISTERS_reg_10_57_inst : DFF_X1 port map( D => n3857, CK => n863, Q => 
                           REGISTERS_10_57_port, QN => n_1650);
   REGISTERS_reg_10_56_inst : DFF_X1 port map( D => n3856, CK => n863, Q => 
                           REGISTERS_10_56_port, QN => n_1651);
   REGISTERS_reg_10_55_inst : DFF_X1 port map( D => n3855, CK => n863, Q => 
                           REGISTERS_10_55_port, QN => n_1652);
   REGISTERS_reg_10_54_inst : DFF_X1 port map( D => n3854, CK => n863, Q => 
                           REGISTERS_10_54_port, QN => n_1653);
   REGISTERS_reg_10_53_inst : DFF_X1 port map( D => n3853, CK => n863, Q => 
                           REGISTERS_10_53_port, QN => n_1654);
   REGISTERS_reg_10_52_inst : DFF_X1 port map( D => n3852, CK => n863, Q => 
                           REGISTERS_10_52_port, QN => n_1655);
   REGISTERS_reg_10_51_inst : DFF_X1 port map( D => n3851, CK => n864, Q => 
                           REGISTERS_10_51_port, QN => n_1656);
   REGISTERS_reg_10_50_inst : DFF_X1 port map( D => n3850, CK => n864, Q => 
                           REGISTERS_10_50_port, QN => n_1657);
   REGISTERS_reg_10_49_inst : DFF_X1 port map( D => n3849, CK => n864, Q => 
                           REGISTERS_10_49_port, QN => n_1658);
   REGISTERS_reg_10_48_inst : DFF_X1 port map( D => n3848, CK => n864, Q => 
                           REGISTERS_10_48_port, QN => n_1659);
   REGISTERS_reg_10_47_inst : DFF_X1 port map( D => n3847, CK => n864, Q => 
                           REGISTERS_10_47_port, QN => n_1660);
   REGISTERS_reg_10_46_inst : DFF_X1 port map( D => n3846, CK => n864, Q => 
                           REGISTERS_10_46_port, QN => n_1661);
   REGISTERS_reg_10_45_inst : DFF_X1 port map( D => n3845, CK => n864, Q => 
                           REGISTERS_10_45_port, QN => n_1662);
   REGISTERS_reg_10_44_inst : DFF_X1 port map( D => n3844, CK => n864, Q => 
                           REGISTERS_10_44_port, QN => n_1663);
   REGISTERS_reg_10_43_inst : DFF_X1 port map( D => n3843, CK => n864, Q => 
                           REGISTERS_10_43_port, QN => n_1664);
   REGISTERS_reg_10_42_inst : DFF_X1 port map( D => n3842, CK => n864, Q => 
                           REGISTERS_10_42_port, QN => n_1665);
   REGISTERS_reg_10_41_inst : DFF_X1 port map( D => n3841, CK => n864, Q => 
                           REGISTERS_10_41_port, QN => n_1666);
   REGISTERS_reg_10_40_inst : DFF_X1 port map( D => n3840, CK => n865, Q => 
                           REGISTERS_10_40_port, QN => n_1667);
   REGISTERS_reg_10_39_inst : DFF_X1 port map( D => n3839, CK => n865, Q => 
                           REGISTERS_10_39_port, QN => n_1668);
   REGISTERS_reg_10_38_inst : DFF_X1 port map( D => n3838, CK => n865, Q => 
                           REGISTERS_10_38_port, QN => n_1669);
   REGISTERS_reg_10_37_inst : DFF_X1 port map( D => n3837, CK => n865, Q => 
                           REGISTERS_10_37_port, QN => n_1670);
   REGISTERS_reg_10_36_inst : DFF_X1 port map( D => n3836, CK => n865, Q => 
                           REGISTERS_10_36_port, QN => n_1671);
   REGISTERS_reg_10_35_inst : DFF_X1 port map( D => n3835, CK => n865, Q => 
                           REGISTERS_10_35_port, QN => n_1672);
   REGISTERS_reg_10_34_inst : DFF_X1 port map( D => n3834, CK => n865, Q => 
                           REGISTERS_10_34_port, QN => n_1673);
   REGISTERS_reg_10_33_inst : DFF_X1 port map( D => n3833, CK => n865, Q => 
                           REGISTERS_10_33_port, QN => n_1674);
   REGISTERS_reg_10_32_inst : DFF_X1 port map( D => n3832, CK => n865, Q => 
                           REGISTERS_10_32_port, QN => n_1675);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n3831, CK => n865, Q => 
                           REGISTERS_10_31_port, QN => n_1676);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n3830, CK => n865, Q => 
                           REGISTERS_10_30_port, QN => n_1677);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n3829, CK => n866, Q => 
                           REGISTERS_10_29_port, QN => n_1678);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n3828, CK => n866, Q => 
                           REGISTERS_10_28_port, QN => n_1679);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n3827, CK => n866, Q => 
                           REGISTERS_10_27_port, QN => n_1680);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n3826, CK => n866, Q => 
                           REGISTERS_10_26_port, QN => n_1681);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n3825, CK => n866, Q => 
                           REGISTERS_10_25_port, QN => n_1682);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n3824, CK => n866, Q => 
                           REGISTERS_10_24_port, QN => n_1683);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n3823, CK => n866, Q => 
                           REGISTERS_10_23_port, QN => n_1684);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n3822, CK => n866, Q => 
                           REGISTERS_10_22_port, QN => n_1685);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n3821, CK => n866, Q => 
                           REGISTERS_10_21_port, QN => n_1686);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n3820, CK => n866, Q => 
                           REGISTERS_10_20_port, QN => n_1687);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n3819, CK => n866, Q => 
                           REGISTERS_10_19_port, QN => n_1688);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n3818, CK => n867, Q => 
                           REGISTERS_10_18_port, QN => n_1689);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n3817, CK => n867, Q => 
                           REGISTERS_10_17_port, QN => n_1690);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n3816, CK => n867, Q => 
                           REGISTERS_10_16_port, QN => n_1691);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n3815, CK => n867, Q => 
                           REGISTERS_10_15_port, QN => n_1692);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n3814, CK => n867, Q => 
                           REGISTERS_10_14_port, QN => n_1693);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n3813, CK => n867, Q => 
                           REGISTERS_10_13_port, QN => n_1694);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n3812, CK => n867, Q => 
                           REGISTERS_10_12_port, QN => n_1695);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n3811, CK => n867, Q => 
                           REGISTERS_10_11_port, QN => n_1696);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n3810, CK => n867, Q => 
                           REGISTERS_10_10_port, QN => n_1697);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n3809, CK => n867, Q => 
                           REGISTERS_10_9_port, QN => n_1698);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n3808, CK => n867, Q => 
                           REGISTERS_10_8_port, QN => n_1699);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n3807, CK => n868, Q => 
                           REGISTERS_10_7_port, QN => n_1700);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n3806, CK => n868, Q => 
                           REGISTERS_10_6_port, QN => n_1701);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n3805, CK => n868, Q => 
                           REGISTERS_10_5_port, QN => n_1702);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n3804, CK => n868, Q => 
                           REGISTERS_10_4_port, QN => n_1703);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n3803, CK => n868, Q => 
                           REGISTERS_10_3_port, QN => n_1704);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n3802, CK => n868, Q => 
                           REGISTERS_10_2_port, QN => n_1705);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n3801, CK => n868, Q => 
                           REGISTERS_10_1_port, QN => n_1706);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n3800, CK => n868, Q => 
                           REGISTERS_10_0_port, QN => n_1707);
   REGISTERS_reg_11_63_inst : DFF_X1 port map( D => n3799, CK => n868, Q => 
                           REGISTERS_11_63_port, QN => n_1708);
   REGISTERS_reg_11_62_inst : DFF_X1 port map( D => n3798, CK => n868, Q => 
                           REGISTERS_11_62_port, QN => n_1709);
   REGISTERS_reg_11_61_inst : DFF_X1 port map( D => n3797, CK => n868, Q => 
                           REGISTERS_11_61_port, QN => n_1710);
   REGISTERS_reg_11_60_inst : DFF_X1 port map( D => n3796, CK => n869, Q => 
                           REGISTERS_11_60_port, QN => n_1711);
   REGISTERS_reg_11_59_inst : DFF_X1 port map( D => n3795, CK => n869, Q => 
                           REGISTERS_11_59_port, QN => n_1712);
   REGISTERS_reg_11_58_inst : DFF_X1 port map( D => n3794, CK => n869, Q => 
                           REGISTERS_11_58_port, QN => n_1713);
   REGISTERS_reg_11_57_inst : DFF_X1 port map( D => n3793, CK => n869, Q => 
                           REGISTERS_11_57_port, QN => n_1714);
   REGISTERS_reg_11_56_inst : DFF_X1 port map( D => n3792, CK => n869, Q => 
                           REGISTERS_11_56_port, QN => n_1715);
   REGISTERS_reg_11_55_inst : DFF_X1 port map( D => n3791, CK => n869, Q => 
                           REGISTERS_11_55_port, QN => n_1716);
   REGISTERS_reg_11_54_inst : DFF_X1 port map( D => n3790, CK => n869, Q => 
                           REGISTERS_11_54_port, QN => n_1717);
   REGISTERS_reg_11_53_inst : DFF_X1 port map( D => n3789, CK => n869, Q => 
                           REGISTERS_11_53_port, QN => n_1718);
   REGISTERS_reg_11_52_inst : DFF_X1 port map( D => n3788, CK => n869, Q => 
                           REGISTERS_11_52_port, QN => n_1719);
   REGISTERS_reg_11_51_inst : DFF_X1 port map( D => n3787, CK => n869, Q => 
                           REGISTERS_11_51_port, QN => n_1720);
   REGISTERS_reg_11_50_inst : DFF_X1 port map( D => n3786, CK => n869, Q => 
                           REGISTERS_11_50_port, QN => n_1721);
   REGISTERS_reg_11_49_inst : DFF_X1 port map( D => n3785, CK => n870, Q => 
                           REGISTERS_11_49_port, QN => n_1722);
   REGISTERS_reg_11_48_inst : DFF_X1 port map( D => n3784, CK => n870, Q => 
                           REGISTERS_11_48_port, QN => n_1723);
   REGISTERS_reg_11_47_inst : DFF_X1 port map( D => n3783, CK => n870, Q => 
                           REGISTERS_11_47_port, QN => n_1724);
   REGISTERS_reg_11_46_inst : DFF_X1 port map( D => n3782, CK => n870, Q => 
                           REGISTERS_11_46_port, QN => n_1725);
   REGISTERS_reg_11_45_inst : DFF_X1 port map( D => n3781, CK => n870, Q => 
                           REGISTERS_11_45_port, QN => n_1726);
   REGISTERS_reg_11_44_inst : DFF_X1 port map( D => n3780, CK => n870, Q => 
                           REGISTERS_11_44_port, QN => n_1727);
   REGISTERS_reg_11_43_inst : DFF_X1 port map( D => n3779, CK => n870, Q => 
                           REGISTERS_11_43_port, QN => n_1728);
   REGISTERS_reg_11_42_inst : DFF_X1 port map( D => n3778, CK => n870, Q => 
                           REGISTERS_11_42_port, QN => n_1729);
   REGISTERS_reg_11_41_inst : DFF_X1 port map( D => n3777, CK => n870, Q => 
                           REGISTERS_11_41_port, QN => n_1730);
   REGISTERS_reg_11_40_inst : DFF_X1 port map( D => n3776, CK => n870, Q => 
                           REGISTERS_11_40_port, QN => n_1731);
   REGISTERS_reg_11_39_inst : DFF_X1 port map( D => n3775, CK => n870, Q => 
                           REGISTERS_11_39_port, QN => n_1732);
   REGISTERS_reg_11_38_inst : DFF_X1 port map( D => n3774, CK => n871, Q => 
                           REGISTERS_11_38_port, QN => n_1733);
   REGISTERS_reg_11_37_inst : DFF_X1 port map( D => n3773, CK => n871, Q => 
                           REGISTERS_11_37_port, QN => n_1734);
   REGISTERS_reg_11_36_inst : DFF_X1 port map( D => n3772, CK => n871, Q => 
                           REGISTERS_11_36_port, QN => n_1735);
   REGISTERS_reg_11_35_inst : DFF_X1 port map( D => n3771, CK => n871, Q => 
                           REGISTERS_11_35_port, QN => n_1736);
   REGISTERS_reg_11_34_inst : DFF_X1 port map( D => n3770, CK => n871, Q => 
                           REGISTERS_11_34_port, QN => n_1737);
   REGISTERS_reg_11_33_inst : DFF_X1 port map( D => n3769, CK => n871, Q => 
                           REGISTERS_11_33_port, QN => n_1738);
   REGISTERS_reg_11_32_inst : DFF_X1 port map( D => n3768, CK => n871, Q => 
                           REGISTERS_11_32_port, QN => n_1739);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n3767, CK => n871, Q => 
                           REGISTERS_11_31_port, QN => n_1740);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n3766, CK => n871, Q => 
                           REGISTERS_11_30_port, QN => n_1741);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n3765, CK => n871, Q => 
                           REGISTERS_11_29_port, QN => n_1742);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n3764, CK => n871, Q => 
                           REGISTERS_11_28_port, QN => n_1743);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n3763, CK => n872, Q => 
                           REGISTERS_11_27_port, QN => n_1744);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n3762, CK => n872, Q => 
                           REGISTERS_11_26_port, QN => n_1745);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n3761, CK => n872, Q => 
                           REGISTERS_11_25_port, QN => n_1746);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n3760, CK => n872, Q => 
                           REGISTERS_11_24_port, QN => n_1747);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n3759, CK => n872, Q => 
                           REGISTERS_11_23_port, QN => n_1748);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n3758, CK => n872, Q => 
                           REGISTERS_11_22_port, QN => n_1749);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n3757, CK => n872, Q => 
                           REGISTERS_11_21_port, QN => n_1750);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n3756, CK => n872, Q => 
                           REGISTERS_11_20_port, QN => n_1751);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n3755, CK => n872, Q => 
                           REGISTERS_11_19_port, QN => n_1752);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n3754, CK => n872, Q => 
                           REGISTERS_11_18_port, QN => n_1753);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n3753, CK => n872, Q => 
                           REGISTERS_11_17_port, QN => n_1754);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n3752, CK => n873, Q => 
                           REGISTERS_11_16_port, QN => n_1755);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n3751, CK => n873, Q => 
                           REGISTERS_11_15_port, QN => n_1756);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n3750, CK => n873, Q => 
                           REGISTERS_11_14_port, QN => n_1757);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n3749, CK => n873, Q => 
                           REGISTERS_11_13_port, QN => n_1758);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n3748, CK => n873, Q => 
                           REGISTERS_11_12_port, QN => n_1759);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n3747, CK => n873, Q => 
                           REGISTERS_11_11_port, QN => n_1760);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n3746, CK => n873, Q => 
                           REGISTERS_11_10_port, QN => n_1761);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n3745, CK => n873, Q => 
                           REGISTERS_11_9_port, QN => n_1762);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n3744, CK => n873, Q => 
                           REGISTERS_11_8_port, QN => n_1763);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n3743, CK => n873, Q => 
                           REGISTERS_11_7_port, QN => n_1764);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n3742, CK => n873, Q => 
                           REGISTERS_11_6_port, QN => n_1765);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n3741, CK => n874, Q => 
                           REGISTERS_11_5_port, QN => n_1766);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n3740, CK => n874, Q => 
                           REGISTERS_11_4_port, QN => n_1767);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n3739, CK => n874, Q => 
                           REGISTERS_11_3_port, QN => n_1768);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n3738, CK => n874, Q => 
                           REGISTERS_11_2_port, QN => n_1769);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n3737, CK => n874, Q => 
                           REGISTERS_11_1_port, QN => n_1770);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n3736, CK => n874, Q => 
                           REGISTERS_11_0_port, QN => n_1771);
   REGISTERS_reg_12_63_inst : DFF_X1 port map( D => n3735, CK => n874, Q => 
                           REGISTERS_12_63_port, QN => n_1772);
   REGISTERS_reg_12_62_inst : DFF_X1 port map( D => n3734, CK => n874, Q => 
                           REGISTERS_12_62_port, QN => n_1773);
   REGISTERS_reg_12_61_inst : DFF_X1 port map( D => n3733, CK => n874, Q => 
                           REGISTERS_12_61_port, QN => n_1774);
   REGISTERS_reg_12_60_inst : DFF_X1 port map( D => n3732, CK => n874, Q => 
                           REGISTERS_12_60_port, QN => n_1775);
   REGISTERS_reg_12_59_inst : DFF_X1 port map( D => n3731, CK => n874, Q => 
                           REGISTERS_12_59_port, QN => n_1776);
   REGISTERS_reg_12_58_inst : DFF_X1 port map( D => n3730, CK => n875, Q => 
                           REGISTERS_12_58_port, QN => n_1777);
   REGISTERS_reg_12_57_inst : DFF_X1 port map( D => n3729, CK => n875, Q => 
                           REGISTERS_12_57_port, QN => n_1778);
   REGISTERS_reg_12_56_inst : DFF_X1 port map( D => n3728, CK => n875, Q => 
                           REGISTERS_12_56_port, QN => n_1779);
   REGISTERS_reg_12_55_inst : DFF_X1 port map( D => n3727, CK => n875, Q => 
                           REGISTERS_12_55_port, QN => n_1780);
   REGISTERS_reg_12_54_inst : DFF_X1 port map( D => n3726, CK => n875, Q => 
                           REGISTERS_12_54_port, QN => n_1781);
   REGISTERS_reg_12_53_inst : DFF_X1 port map( D => n3725, CK => n875, Q => 
                           REGISTERS_12_53_port, QN => n_1782);
   REGISTERS_reg_12_52_inst : DFF_X1 port map( D => n3724, CK => n875, Q => 
                           REGISTERS_12_52_port, QN => n_1783);
   REGISTERS_reg_12_51_inst : DFF_X1 port map( D => n3723, CK => n875, Q => 
                           REGISTERS_12_51_port, QN => n_1784);
   REGISTERS_reg_12_50_inst : DFF_X1 port map( D => n3722, CK => n875, Q => 
                           REGISTERS_12_50_port, QN => n_1785);
   REGISTERS_reg_12_49_inst : DFF_X1 port map( D => n3721, CK => n875, Q => 
                           REGISTERS_12_49_port, QN => n_1786);
   REGISTERS_reg_12_48_inst : DFF_X1 port map( D => n3720, CK => n875, Q => 
                           REGISTERS_12_48_port, QN => n_1787);
   REGISTERS_reg_12_47_inst : DFF_X1 port map( D => n3719, CK => n876, Q => 
                           REGISTERS_12_47_port, QN => n_1788);
   REGISTERS_reg_12_46_inst : DFF_X1 port map( D => n3718, CK => n876, Q => 
                           REGISTERS_12_46_port, QN => n_1789);
   REGISTERS_reg_12_45_inst : DFF_X1 port map( D => n3717, CK => n876, Q => 
                           REGISTERS_12_45_port, QN => n_1790);
   REGISTERS_reg_12_44_inst : DFF_X1 port map( D => n3716, CK => n876, Q => 
                           REGISTERS_12_44_port, QN => n_1791);
   REGISTERS_reg_12_43_inst : DFF_X1 port map( D => n3715, CK => n876, Q => 
                           REGISTERS_12_43_port, QN => n_1792);
   REGISTERS_reg_12_42_inst : DFF_X1 port map( D => n3714, CK => n876, Q => 
                           REGISTERS_12_42_port, QN => n_1793);
   REGISTERS_reg_12_41_inst : DFF_X1 port map( D => n3713, CK => n876, Q => 
                           REGISTERS_12_41_port, QN => n_1794);
   REGISTERS_reg_12_40_inst : DFF_X1 port map( D => n3712, CK => n876, Q => 
                           REGISTERS_12_40_port, QN => n_1795);
   REGISTERS_reg_12_39_inst : DFF_X1 port map( D => n3711, CK => n876, Q => 
                           REGISTERS_12_39_port, QN => n_1796);
   REGISTERS_reg_12_38_inst : DFF_X1 port map( D => n3710, CK => n876, Q => 
                           REGISTERS_12_38_port, QN => n_1797);
   REGISTERS_reg_12_37_inst : DFF_X1 port map( D => n3709, CK => n876, Q => 
                           REGISTERS_12_37_port, QN => n_1798);
   REGISTERS_reg_12_36_inst : DFF_X1 port map( D => n3708, CK => n877, Q => 
                           REGISTERS_12_36_port, QN => n_1799);
   REGISTERS_reg_12_35_inst : DFF_X1 port map( D => n3707, CK => n877, Q => 
                           REGISTERS_12_35_port, QN => n_1800);
   REGISTERS_reg_12_34_inst : DFF_X1 port map( D => n3706, CK => n877, Q => 
                           REGISTERS_12_34_port, QN => n_1801);
   REGISTERS_reg_12_33_inst : DFF_X1 port map( D => n3705, CK => n877, Q => 
                           REGISTERS_12_33_port, QN => n_1802);
   REGISTERS_reg_12_32_inst : DFF_X1 port map( D => n3704, CK => n877, Q => 
                           REGISTERS_12_32_port, QN => n_1803);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n3703, CK => n877, Q => 
                           REGISTERS_12_31_port, QN => n_1804);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n3702, CK => n877, Q => 
                           REGISTERS_12_30_port, QN => n_1805);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n3701, CK => n877, Q => 
                           REGISTERS_12_29_port, QN => n_1806);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n3700, CK => n877, Q => 
                           REGISTERS_12_28_port, QN => n_1807);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n3699, CK => n877, Q => 
                           REGISTERS_12_27_port, QN => n_1808);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n3698, CK => n877, Q => 
                           REGISTERS_12_26_port, QN => n_1809);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n3697, CK => n878, Q => 
                           REGISTERS_12_25_port, QN => n_1810);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n3696, CK => n878, Q => 
                           REGISTERS_12_24_port, QN => n_1811);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n3695, CK => n878, Q => 
                           REGISTERS_12_23_port, QN => n_1812);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n3694, CK => n878, Q => 
                           REGISTERS_12_22_port, QN => n_1813);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n3693, CK => n878, Q => 
                           REGISTERS_12_21_port, QN => n_1814);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n3692, CK => n878, Q => 
                           REGISTERS_12_20_port, QN => n_1815);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n3691, CK => n878, Q => 
                           REGISTERS_12_19_port, QN => n_1816);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n3690, CK => n878, Q => 
                           REGISTERS_12_18_port, QN => n_1817);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n3689, CK => n878, Q => 
                           REGISTERS_12_17_port, QN => n_1818);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n3688, CK => n878, Q => 
                           REGISTERS_12_16_port, QN => n_1819);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n3687, CK => n878, Q => 
                           REGISTERS_12_15_port, QN => n_1820);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n3686, CK => n879, Q => 
                           REGISTERS_12_14_port, QN => n_1821);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n3685, CK => n879, Q => 
                           REGISTERS_12_13_port, QN => n_1822);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n3684, CK => n879, Q => 
                           REGISTERS_12_12_port, QN => n_1823);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n3683, CK => n879, Q => 
                           REGISTERS_12_11_port, QN => n_1824);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n3682, CK => n879, Q => 
                           REGISTERS_12_10_port, QN => n_1825);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n3681, CK => n879, Q => 
                           REGISTERS_12_9_port, QN => n_1826);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n3680, CK => n879, Q => 
                           REGISTERS_12_8_port, QN => n_1827);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n3679, CK => n879, Q => 
                           REGISTERS_12_7_port, QN => n_1828);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n3678, CK => n879, Q => 
                           REGISTERS_12_6_port, QN => n_1829);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n3677, CK => n879, Q => 
                           REGISTERS_12_5_port, QN => n_1830);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n3676, CK => n879, Q => 
                           REGISTERS_12_4_port, QN => n_1831);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n3675, CK => n880, Q => 
                           REGISTERS_12_3_port, QN => n_1832);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n3674, CK => n880, Q => 
                           REGISTERS_12_2_port, QN => n_1833);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n3673, CK => n880, Q => 
                           REGISTERS_12_1_port, QN => n_1834);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n3672, CK => n880, Q => 
                           REGISTERS_12_0_port, QN => n_1835);
   REGISTERS_reg_13_63_inst : DFF_X1 port map( D => n3671, CK => n880, Q => 
                           REGISTERS_13_63_port, QN => n_1836);
   REGISTERS_reg_13_62_inst : DFF_X1 port map( D => n3670, CK => n880, Q => 
                           REGISTERS_13_62_port, QN => n_1837);
   REGISTERS_reg_13_61_inst : DFF_X1 port map( D => n3669, CK => n880, Q => 
                           REGISTERS_13_61_port, QN => n_1838);
   REGISTERS_reg_13_60_inst : DFF_X1 port map( D => n3668, CK => n880, Q => 
                           REGISTERS_13_60_port, QN => n_1839);
   REGISTERS_reg_13_59_inst : DFF_X1 port map( D => n3667, CK => n880, Q => 
                           REGISTERS_13_59_port, QN => n_1840);
   REGISTERS_reg_13_58_inst : DFF_X1 port map( D => n3666, CK => n880, Q => 
                           REGISTERS_13_58_port, QN => n_1841);
   REGISTERS_reg_13_57_inst : DFF_X1 port map( D => n3665, CK => n880, Q => 
                           REGISTERS_13_57_port, QN => n_1842);
   REGISTERS_reg_13_56_inst : DFF_X1 port map( D => n3664, CK => n881, Q => 
                           REGISTERS_13_56_port, QN => n_1843);
   REGISTERS_reg_13_55_inst : DFF_X1 port map( D => n3663, CK => n881, Q => 
                           REGISTERS_13_55_port, QN => n_1844);
   REGISTERS_reg_13_54_inst : DFF_X1 port map( D => n3662, CK => n881, Q => 
                           REGISTERS_13_54_port, QN => n_1845);
   REGISTERS_reg_13_53_inst : DFF_X1 port map( D => n3661, CK => n881, Q => 
                           REGISTERS_13_53_port, QN => n_1846);
   REGISTERS_reg_13_52_inst : DFF_X1 port map( D => n3660, CK => n881, Q => 
                           REGISTERS_13_52_port, QN => n_1847);
   REGISTERS_reg_13_51_inst : DFF_X1 port map( D => n3659, CK => n881, Q => 
                           REGISTERS_13_51_port, QN => n_1848);
   REGISTERS_reg_13_50_inst : DFF_X1 port map( D => n3658, CK => n881, Q => 
                           REGISTERS_13_50_port, QN => n_1849);
   REGISTERS_reg_13_49_inst : DFF_X1 port map( D => n3657, CK => n881, Q => 
                           REGISTERS_13_49_port, QN => n_1850);
   REGISTERS_reg_13_48_inst : DFF_X1 port map( D => n3656, CK => n881, Q => 
                           REGISTERS_13_48_port, QN => n_1851);
   REGISTERS_reg_13_47_inst : DFF_X1 port map( D => n3655, CK => n881, Q => 
                           REGISTERS_13_47_port, QN => n_1852);
   REGISTERS_reg_13_46_inst : DFF_X1 port map( D => n3654, CK => n881, Q => 
                           REGISTERS_13_46_port, QN => n_1853);
   REGISTERS_reg_13_45_inst : DFF_X1 port map( D => n3653, CK => n882, Q => 
                           REGISTERS_13_45_port, QN => n_1854);
   REGISTERS_reg_13_44_inst : DFF_X1 port map( D => n3652, CK => n882, Q => 
                           REGISTERS_13_44_port, QN => n_1855);
   REGISTERS_reg_13_43_inst : DFF_X1 port map( D => n3651, CK => n882, Q => 
                           REGISTERS_13_43_port, QN => n_1856);
   REGISTERS_reg_13_42_inst : DFF_X1 port map( D => n3650, CK => n882, Q => 
                           REGISTERS_13_42_port, QN => n_1857);
   REGISTERS_reg_13_41_inst : DFF_X1 port map( D => n3649, CK => n882, Q => 
                           REGISTERS_13_41_port, QN => n_1858);
   REGISTERS_reg_13_40_inst : DFF_X1 port map( D => n3648, CK => n882, Q => 
                           REGISTERS_13_40_port, QN => n_1859);
   REGISTERS_reg_13_39_inst : DFF_X1 port map( D => n3647, CK => n882, Q => 
                           REGISTERS_13_39_port, QN => n_1860);
   REGISTERS_reg_13_38_inst : DFF_X1 port map( D => n3646, CK => n882, Q => 
                           REGISTERS_13_38_port, QN => n_1861);
   REGISTERS_reg_13_37_inst : DFF_X1 port map( D => n3645, CK => n882, Q => 
                           REGISTERS_13_37_port, QN => n_1862);
   REGISTERS_reg_13_36_inst : DFF_X1 port map( D => n3644, CK => n882, Q => 
                           REGISTERS_13_36_port, QN => n_1863);
   REGISTERS_reg_13_35_inst : DFF_X1 port map( D => n3643, CK => n882, Q => 
                           REGISTERS_13_35_port, QN => n_1864);
   REGISTERS_reg_13_34_inst : DFF_X1 port map( D => n3642, CK => n883, Q => 
                           REGISTERS_13_34_port, QN => n_1865);
   REGISTERS_reg_13_33_inst : DFF_X1 port map( D => n3641, CK => n883, Q => 
                           REGISTERS_13_33_port, QN => n_1866);
   REGISTERS_reg_13_32_inst : DFF_X1 port map( D => n3640, CK => n883, Q => 
                           REGISTERS_13_32_port, QN => n_1867);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n3639, CK => n883, Q => 
                           REGISTERS_13_31_port, QN => n_1868);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n3638, CK => n883, Q => 
                           REGISTERS_13_30_port, QN => n_1869);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n3637, CK => n883, Q => 
                           REGISTERS_13_29_port, QN => n_1870);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n3636, CK => n883, Q => 
                           REGISTERS_13_28_port, QN => n_1871);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n3635, CK => n883, Q => 
                           REGISTERS_13_27_port, QN => n_1872);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n3634, CK => n883, Q => 
                           REGISTERS_13_26_port, QN => n_1873);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n3633, CK => n883, Q => 
                           REGISTERS_13_25_port, QN => n_1874);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n3632, CK => n883, Q => 
                           REGISTERS_13_24_port, QN => n_1875);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n3631, CK => n884, Q => 
                           REGISTERS_13_23_port, QN => n_1876);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n3630, CK => n884, Q => 
                           REGISTERS_13_22_port, QN => n_1877);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n3629, CK => n884, Q => 
                           REGISTERS_13_21_port, QN => n_1878);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n3628, CK => n884, Q => 
                           REGISTERS_13_20_port, QN => n_1879);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n3627, CK => n884, Q => 
                           REGISTERS_13_19_port, QN => n_1880);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n3626, CK => n884, Q => 
                           REGISTERS_13_18_port, QN => n_1881);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n3625, CK => n884, Q => 
                           REGISTERS_13_17_port, QN => n_1882);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n3624, CK => n884, Q => 
                           REGISTERS_13_16_port, QN => n_1883);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n3623, CK => n884, Q => 
                           REGISTERS_13_15_port, QN => n_1884);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n3622, CK => n884, Q => 
                           REGISTERS_13_14_port, QN => n_1885);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n3621, CK => n884, Q => 
                           REGISTERS_13_13_port, QN => n_1886);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n3620, CK => n885, Q => 
                           REGISTERS_13_12_port, QN => n_1887);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n3619, CK => n885, Q => 
                           REGISTERS_13_11_port, QN => n_1888);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n3618, CK => n885, Q => 
                           REGISTERS_13_10_port, QN => n_1889);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n3617, CK => n885, Q => 
                           REGISTERS_13_9_port, QN => n_1890);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n3616, CK => n885, Q => 
                           REGISTERS_13_8_port, QN => n_1891);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n3615, CK => n885, Q => 
                           REGISTERS_13_7_port, QN => n_1892);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n3614, CK => n885, Q => 
                           REGISTERS_13_6_port, QN => n_1893);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n3613, CK => n885, Q => 
                           REGISTERS_13_5_port, QN => n_1894);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n3612, CK => n885, Q => 
                           REGISTERS_13_4_port, QN => n_1895);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n3611, CK => n885, Q => 
                           REGISTERS_13_3_port, QN => n_1896);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n3610, CK => n885, Q => 
                           REGISTERS_13_2_port, QN => n_1897);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n3609, CK => n886, Q => 
                           REGISTERS_13_1_port, QN => n_1898);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n3608, CK => n886, Q => 
                           REGISTERS_13_0_port, QN => n_1899);
   REGISTERS_reg_14_63_inst : DFF_X1 port map( D => n3607, CK => n886, Q => 
                           REGISTERS_14_63_port, QN => n_1900);
   REGISTERS_reg_14_62_inst : DFF_X1 port map( D => n3606, CK => n886, Q => 
                           REGISTERS_14_62_port, QN => n_1901);
   REGISTERS_reg_14_61_inst : DFF_X1 port map( D => n3605, CK => n886, Q => 
                           REGISTERS_14_61_port, QN => n_1902);
   REGISTERS_reg_14_60_inst : DFF_X1 port map( D => n3604, CK => n886, Q => 
                           REGISTERS_14_60_port, QN => n_1903);
   REGISTERS_reg_14_59_inst : DFF_X1 port map( D => n3603, CK => n886, Q => 
                           REGISTERS_14_59_port, QN => n_1904);
   REGISTERS_reg_14_58_inst : DFF_X1 port map( D => n3602, CK => n886, Q => 
                           REGISTERS_14_58_port, QN => n_1905);
   REGISTERS_reg_14_57_inst : DFF_X1 port map( D => n3601, CK => n886, Q => 
                           REGISTERS_14_57_port, QN => n_1906);
   REGISTERS_reg_14_56_inst : DFF_X1 port map( D => n3600, CK => n886, Q => 
                           REGISTERS_14_56_port, QN => n_1907);
   REGISTERS_reg_14_55_inst : DFF_X1 port map( D => n3599, CK => n886, Q => 
                           REGISTERS_14_55_port, QN => n_1908);
   REGISTERS_reg_14_54_inst : DFF_X1 port map( D => n3598, CK => n887, Q => 
                           REGISTERS_14_54_port, QN => n_1909);
   REGISTERS_reg_14_53_inst : DFF_X1 port map( D => n3597, CK => n887, Q => 
                           REGISTERS_14_53_port, QN => n_1910);
   REGISTERS_reg_14_52_inst : DFF_X1 port map( D => n3596, CK => n887, Q => 
                           REGISTERS_14_52_port, QN => n_1911);
   REGISTERS_reg_14_51_inst : DFF_X1 port map( D => n3595, CK => n887, Q => 
                           REGISTERS_14_51_port, QN => n_1912);
   REGISTERS_reg_14_50_inst : DFF_X1 port map( D => n3594, CK => n887, Q => 
                           REGISTERS_14_50_port, QN => n_1913);
   REGISTERS_reg_14_49_inst : DFF_X1 port map( D => n3593, CK => n887, Q => 
                           REGISTERS_14_49_port, QN => n_1914);
   REGISTERS_reg_14_48_inst : DFF_X1 port map( D => n3592, CK => n887, Q => 
                           REGISTERS_14_48_port, QN => n_1915);
   REGISTERS_reg_14_47_inst : DFF_X1 port map( D => n3591, CK => n887, Q => 
                           REGISTERS_14_47_port, QN => n_1916);
   REGISTERS_reg_14_46_inst : DFF_X1 port map( D => n3590, CK => n887, Q => 
                           REGISTERS_14_46_port, QN => n_1917);
   REGISTERS_reg_14_45_inst : DFF_X1 port map( D => n3589, CK => n887, Q => 
                           REGISTERS_14_45_port, QN => n_1918);
   REGISTERS_reg_14_44_inst : DFF_X1 port map( D => n3588, CK => n887, Q => 
                           REGISTERS_14_44_port, QN => n_1919);
   REGISTERS_reg_14_43_inst : DFF_X1 port map( D => n3587, CK => n888, Q => 
                           REGISTERS_14_43_port, QN => n_1920);
   REGISTERS_reg_14_42_inst : DFF_X1 port map( D => n3586, CK => n888, Q => 
                           REGISTERS_14_42_port, QN => n_1921);
   REGISTERS_reg_14_41_inst : DFF_X1 port map( D => n3585, CK => n888, Q => 
                           REGISTERS_14_41_port, QN => n_1922);
   REGISTERS_reg_14_40_inst : DFF_X1 port map( D => n3584, CK => n888, Q => 
                           REGISTERS_14_40_port, QN => n_1923);
   REGISTERS_reg_14_39_inst : DFF_X1 port map( D => n3583, CK => n888, Q => 
                           REGISTERS_14_39_port, QN => n_1924);
   REGISTERS_reg_14_38_inst : DFF_X1 port map( D => n3582, CK => n888, Q => 
                           REGISTERS_14_38_port, QN => n_1925);
   REGISTERS_reg_14_37_inst : DFF_X1 port map( D => n3581, CK => n888, Q => 
                           REGISTERS_14_37_port, QN => n_1926);
   REGISTERS_reg_14_36_inst : DFF_X1 port map( D => n3580, CK => n888, Q => 
                           REGISTERS_14_36_port, QN => n_1927);
   REGISTERS_reg_14_35_inst : DFF_X1 port map( D => n3579, CK => n888, Q => 
                           REGISTERS_14_35_port, QN => n_1928);
   REGISTERS_reg_14_34_inst : DFF_X1 port map( D => n3578, CK => n888, Q => 
                           REGISTERS_14_34_port, QN => n_1929);
   REGISTERS_reg_14_33_inst : DFF_X1 port map( D => n3577, CK => n888, Q => 
                           REGISTERS_14_33_port, QN => n_1930);
   REGISTERS_reg_14_32_inst : DFF_X1 port map( D => n3576, CK => n889, Q => 
                           REGISTERS_14_32_port, QN => n_1931);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n3575, CK => n889, Q => 
                           REGISTERS_14_31_port, QN => n_1932);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n3574, CK => n889, Q => 
                           REGISTERS_14_30_port, QN => n_1933);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n3573, CK => n889, Q => 
                           REGISTERS_14_29_port, QN => n_1934);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n3572, CK => n889, Q => 
                           REGISTERS_14_28_port, QN => n_1935);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n3571, CK => n889, Q => 
                           REGISTERS_14_27_port, QN => n_1936);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n3570, CK => n889, Q => 
                           REGISTERS_14_26_port, QN => n_1937);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n3569, CK => n889, Q => 
                           REGISTERS_14_25_port, QN => n_1938);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n3568, CK => n889, Q => 
                           REGISTERS_14_24_port, QN => n_1939);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n3567, CK => n889, Q => 
                           REGISTERS_14_23_port, QN => n_1940);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n3566, CK => n889, Q => 
                           REGISTERS_14_22_port, QN => n_1941);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n3565, CK => n890, Q => 
                           REGISTERS_14_21_port, QN => n_1942);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n3564, CK => n890, Q => 
                           REGISTERS_14_20_port, QN => n_1943);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n3563, CK => n890, Q => 
                           REGISTERS_14_19_port, QN => n_1944);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n3562, CK => n890, Q => 
                           REGISTERS_14_18_port, QN => n_1945);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n3561, CK => n890, Q => 
                           REGISTERS_14_17_port, QN => n_1946);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n3560, CK => n890, Q => 
                           REGISTERS_14_16_port, QN => n_1947);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n3559, CK => n890, Q => 
                           REGISTERS_14_15_port, QN => n_1948);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n3558, CK => n890, Q => 
                           REGISTERS_14_14_port, QN => n_1949);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n3557, CK => n890, Q => 
                           REGISTERS_14_13_port, QN => n_1950);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n3556, CK => n890, Q => 
                           REGISTERS_14_12_port, QN => n_1951);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n3555, CK => n890, Q => 
                           REGISTERS_14_11_port, QN => n_1952);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n3554, CK => n891, Q => 
                           REGISTERS_14_10_port, QN => n_1953);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n3553, CK => n891, Q => 
                           REGISTERS_14_9_port, QN => n_1954);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n3552, CK => n891, Q => 
                           REGISTERS_14_8_port, QN => n_1955);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n3551, CK => n891, Q => 
                           REGISTERS_14_7_port, QN => n_1956);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n3550, CK => n891, Q => 
                           REGISTERS_14_6_port, QN => n_1957);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n3549, CK => n891, Q => 
                           REGISTERS_14_5_port, QN => n_1958);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n3548, CK => n891, Q => 
                           REGISTERS_14_4_port, QN => n_1959);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n3547, CK => n891, Q => 
                           REGISTERS_14_3_port, QN => n_1960);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n3546, CK => n891, Q => 
                           REGISTERS_14_2_port, QN => n_1961);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n3545, CK => n891, Q => 
                           REGISTERS_14_1_port, QN => n_1962);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n3544, CK => n891, Q => 
                           REGISTERS_14_0_port, QN => n_1963);
   REGISTERS_reg_15_63_inst : DFF_X1 port map( D => n3543, CK => n892, Q => 
                           REGISTERS_15_63_port, QN => n_1964);
   REGISTERS_reg_15_62_inst : DFF_X1 port map( D => n3542, CK => n892, Q => 
                           REGISTERS_15_62_port, QN => n_1965);
   REGISTERS_reg_15_61_inst : DFF_X1 port map( D => n3541, CK => n892, Q => 
                           REGISTERS_15_61_port, QN => n_1966);
   REGISTERS_reg_15_60_inst : DFF_X1 port map( D => n3540, CK => n892, Q => 
                           REGISTERS_15_60_port, QN => n_1967);
   REGISTERS_reg_15_59_inst : DFF_X1 port map( D => n3539, CK => n892, Q => 
                           REGISTERS_15_59_port, QN => n_1968);
   REGISTERS_reg_15_58_inst : DFF_X1 port map( D => n3538, CK => n892, Q => 
                           REGISTERS_15_58_port, QN => n_1969);
   REGISTERS_reg_15_57_inst : DFF_X1 port map( D => n3537, CK => n892, Q => 
                           REGISTERS_15_57_port, QN => n_1970);
   REGISTERS_reg_15_56_inst : DFF_X1 port map( D => n3536, CK => n892, Q => 
                           REGISTERS_15_56_port, QN => n_1971);
   REGISTERS_reg_15_55_inst : DFF_X1 port map( D => n3535, CK => n892, Q => 
                           REGISTERS_15_55_port, QN => n_1972);
   REGISTERS_reg_15_54_inst : DFF_X1 port map( D => n3534, CK => n892, Q => 
                           REGISTERS_15_54_port, QN => n_1973);
   REGISTERS_reg_15_53_inst : DFF_X1 port map( D => n3533, CK => n892, Q => 
                           REGISTERS_15_53_port, QN => n_1974);
   REGISTERS_reg_15_52_inst : DFF_X1 port map( D => n3532, CK => n893, Q => 
                           REGISTERS_15_52_port, QN => n_1975);
   REGISTERS_reg_15_51_inst : DFF_X1 port map( D => n3531, CK => n893, Q => 
                           REGISTERS_15_51_port, QN => n_1976);
   REGISTERS_reg_15_50_inst : DFF_X1 port map( D => n3530, CK => n893, Q => 
                           REGISTERS_15_50_port, QN => n_1977);
   REGISTERS_reg_15_49_inst : DFF_X1 port map( D => n3529, CK => n893, Q => 
                           REGISTERS_15_49_port, QN => n_1978);
   REGISTERS_reg_15_48_inst : DFF_X1 port map( D => n3528, CK => n893, Q => 
                           REGISTERS_15_48_port, QN => n_1979);
   REGISTERS_reg_15_47_inst : DFF_X1 port map( D => n3527, CK => n893, Q => 
                           REGISTERS_15_47_port, QN => n_1980);
   REGISTERS_reg_15_46_inst : DFF_X1 port map( D => n3526, CK => n893, Q => 
                           REGISTERS_15_46_port, QN => n_1981);
   REGISTERS_reg_15_45_inst : DFF_X1 port map( D => n3525, CK => n893, Q => 
                           REGISTERS_15_45_port, QN => n_1982);
   REGISTERS_reg_15_44_inst : DFF_X1 port map( D => n3524, CK => n893, Q => 
                           REGISTERS_15_44_port, QN => n_1983);
   REGISTERS_reg_15_43_inst : DFF_X1 port map( D => n3523, CK => n893, Q => 
                           REGISTERS_15_43_port, QN => n_1984);
   REGISTERS_reg_15_42_inst : DFF_X1 port map( D => n3522, CK => n893, Q => 
                           REGISTERS_15_42_port, QN => n_1985);
   REGISTERS_reg_15_41_inst : DFF_X1 port map( D => n3521, CK => n894, Q => 
                           REGISTERS_15_41_port, QN => n_1986);
   REGISTERS_reg_15_40_inst : DFF_X1 port map( D => n3520, CK => n894, Q => 
                           REGISTERS_15_40_port, QN => n_1987);
   REGISTERS_reg_15_39_inst : DFF_X1 port map( D => n3519, CK => n894, Q => 
                           REGISTERS_15_39_port, QN => n_1988);
   REGISTERS_reg_15_38_inst : DFF_X1 port map( D => n3518, CK => n894, Q => 
                           REGISTERS_15_38_port, QN => n_1989);
   REGISTERS_reg_15_37_inst : DFF_X1 port map( D => n3517, CK => n894, Q => 
                           REGISTERS_15_37_port, QN => n_1990);
   REGISTERS_reg_15_36_inst : DFF_X1 port map( D => n3516, CK => n894, Q => 
                           REGISTERS_15_36_port, QN => n_1991);
   REGISTERS_reg_15_35_inst : DFF_X1 port map( D => n3515, CK => n894, Q => 
                           REGISTERS_15_35_port, QN => n_1992);
   REGISTERS_reg_15_34_inst : DFF_X1 port map( D => n3514, CK => n894, Q => 
                           REGISTERS_15_34_port, QN => n_1993);
   REGISTERS_reg_15_33_inst : DFF_X1 port map( D => n3513, CK => n894, Q => 
                           REGISTERS_15_33_port, QN => n_1994);
   REGISTERS_reg_15_32_inst : DFF_X1 port map( D => n3512, CK => n894, Q => 
                           REGISTERS_15_32_port, QN => n_1995);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n3511, CK => n894, Q => 
                           REGISTERS_15_31_port, QN => n_1996);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n3510, CK => n895, Q => 
                           REGISTERS_15_30_port, QN => n_1997);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n3509, CK => n895, Q => 
                           REGISTERS_15_29_port, QN => n_1998);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n3508, CK => n895, Q => 
                           REGISTERS_15_28_port, QN => n_1999);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n3507, CK => n895, Q => 
                           REGISTERS_15_27_port, QN => n_2000);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n3506, CK => n895, Q => 
                           REGISTERS_15_26_port, QN => n_2001);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n3505, CK => n895, Q => 
                           REGISTERS_15_25_port, QN => n_2002);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n3504, CK => n895, Q => 
                           REGISTERS_15_24_port, QN => n_2003);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n3503, CK => n895, Q => 
                           REGISTERS_15_23_port, QN => n_2004);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n3502, CK => n895, Q => 
                           REGISTERS_15_22_port, QN => n_2005);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n3501, CK => n895, Q => 
                           REGISTERS_15_21_port, QN => n_2006);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n3500, CK => n895, Q => 
                           REGISTERS_15_20_port, QN => n_2007);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n3499, CK => n896, Q => 
                           REGISTERS_15_19_port, QN => n_2008);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n3498, CK => n896, Q => 
                           REGISTERS_15_18_port, QN => n_2009);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n3497, CK => n896, Q => 
                           REGISTERS_15_17_port, QN => n_2010);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n3496, CK => n896, Q => 
                           REGISTERS_15_16_port, QN => n_2011);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n3495, CK => n896, Q => 
                           REGISTERS_15_15_port, QN => n_2012);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n3494, CK => n896, Q => 
                           REGISTERS_15_14_port, QN => n_2013);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n3493, CK => n896, Q => 
                           REGISTERS_15_13_port, QN => n_2014);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n3492, CK => n896, Q => 
                           REGISTERS_15_12_port, QN => n_2015);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n3491, CK => n896, Q => 
                           REGISTERS_15_11_port, QN => n_2016);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n3490, CK => n896, Q => 
                           REGISTERS_15_10_port, QN => n_2017);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n3489, CK => n896, Q => 
                           REGISTERS_15_9_port, QN => n_2018);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n3488, CK => n897, Q => 
                           REGISTERS_15_8_port, QN => n_2019);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n3487, CK => n897, Q => 
                           REGISTERS_15_7_port, QN => n_2020);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n3486, CK => n897, Q => 
                           REGISTERS_15_6_port, QN => n_2021);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n3485, CK => n897, Q => 
                           REGISTERS_15_5_port, QN => n_2022);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n3484, CK => n897, Q => 
                           REGISTERS_15_4_port, QN => n_2023);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n3483, CK => n897, Q => 
                           REGISTERS_15_3_port, QN => n_2024);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n3482, CK => n897, Q => 
                           REGISTERS_15_2_port, QN => n_2025);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n3481, CK => n897, Q => 
                           REGISTERS_15_1_port, QN => n_2026);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n3480, CK => n897, Q => 
                           REGISTERS_15_0_port, QN => n_2027);
   REGISTERS_reg_16_63_inst : DFF_X1 port map( D => n3479, CK => n758, Q => 
                           REGISTERS_16_63_port, QN => n_2028);
   REGISTERS_reg_16_62_inst : DFF_X1 port map( D => n3478, CK => n758, Q => 
                           REGISTERS_16_62_port, QN => n_2029);
   REGISTERS_reg_16_61_inst : DFF_X1 port map( D => n3477, CK => n758, Q => 
                           REGISTERS_16_61_port, QN => n_2030);
   REGISTERS_reg_16_60_inst : DFF_X1 port map( D => n3476, CK => n758, Q => 
                           REGISTERS_16_60_port, QN => n_2031);
   REGISTERS_reg_16_59_inst : DFF_X1 port map( D => n3475, CK => n758, Q => 
                           REGISTERS_16_59_port, QN => n_2032);
   REGISTERS_reg_16_58_inst : DFF_X1 port map( D => n3474, CK => n758, Q => 
                           REGISTERS_16_58_port, QN => n_2033);
   REGISTERS_reg_16_57_inst : DFF_X1 port map( D => n3473, CK => n758, Q => 
                           REGISTERS_16_57_port, QN => n_2034);
   REGISTERS_reg_16_56_inst : DFF_X1 port map( D => n3472, CK => n758, Q => 
                           REGISTERS_16_56_port, QN => n_2035);
   REGISTERS_reg_16_55_inst : DFF_X1 port map( D => n3471, CK => n758, Q => 
                           REGISTERS_16_55_port, QN => n_2036);
   REGISTERS_reg_16_54_inst : DFF_X1 port map( D => n3470, CK => n759, Q => 
                           REGISTERS_16_54_port, QN => n_2037);
   REGISTERS_reg_16_53_inst : DFF_X1 port map( D => n3469, CK => n759, Q => 
                           REGISTERS_16_53_port, QN => n_2038);
   REGISTERS_reg_16_52_inst : DFF_X1 port map( D => n3468, CK => n759, Q => 
                           REGISTERS_16_52_port, QN => n_2039);
   REGISTERS_reg_16_51_inst : DFF_X1 port map( D => n3467, CK => n759, Q => 
                           REGISTERS_16_51_port, QN => n_2040);
   REGISTERS_reg_16_50_inst : DFF_X1 port map( D => n3466, CK => n759, Q => 
                           REGISTERS_16_50_port, QN => n_2041);
   REGISTERS_reg_16_49_inst : DFF_X1 port map( D => n3465, CK => n759, Q => 
                           REGISTERS_16_49_port, QN => n_2042);
   REGISTERS_reg_16_48_inst : DFF_X1 port map( D => n3464, CK => n759, Q => 
                           REGISTERS_16_48_port, QN => n_2043);
   REGISTERS_reg_16_47_inst : DFF_X1 port map( D => n3463, CK => n759, Q => 
                           REGISTERS_16_47_port, QN => n_2044);
   REGISTERS_reg_16_46_inst : DFF_X1 port map( D => n3462, CK => n759, Q => 
                           REGISTERS_16_46_port, QN => n_2045);
   REGISTERS_reg_16_45_inst : DFF_X1 port map( D => n3461, CK => n759, Q => 
                           REGISTERS_16_45_port, QN => n_2046);
   REGISTERS_reg_16_44_inst : DFF_X1 port map( D => n3460, CK => n759, Q => 
                           REGISTERS_16_44_port, QN => n_2047);
   REGISTERS_reg_16_43_inst : DFF_X1 port map( D => n3459, CK => n760, Q => 
                           REGISTERS_16_43_port, QN => n_2048);
   REGISTERS_reg_16_42_inst : DFF_X1 port map( D => n3458, CK => n760, Q => 
                           REGISTERS_16_42_port, QN => n_2049);
   REGISTERS_reg_16_41_inst : DFF_X1 port map( D => n3457, CK => n760, Q => 
                           REGISTERS_16_41_port, QN => n_2050);
   REGISTERS_reg_16_40_inst : DFF_X1 port map( D => n3456, CK => n760, Q => 
                           REGISTERS_16_40_port, QN => n_2051);
   REGISTERS_reg_16_39_inst : DFF_X1 port map( D => n3455, CK => n760, Q => 
                           REGISTERS_16_39_port, QN => n_2052);
   REGISTERS_reg_16_38_inst : DFF_X1 port map( D => n3454, CK => n760, Q => 
                           REGISTERS_16_38_port, QN => n_2053);
   REGISTERS_reg_16_37_inst : DFF_X1 port map( D => n3453, CK => n760, Q => 
                           REGISTERS_16_37_port, QN => n_2054);
   REGISTERS_reg_16_36_inst : DFF_X1 port map( D => n3452, CK => n760, Q => 
                           REGISTERS_16_36_port, QN => n_2055);
   REGISTERS_reg_16_35_inst : DFF_X1 port map( D => n3451, CK => n760, Q => 
                           REGISTERS_16_35_port, QN => n_2056);
   REGISTERS_reg_16_34_inst : DFF_X1 port map( D => n3450, CK => n760, Q => 
                           REGISTERS_16_34_port, QN => n_2057);
   REGISTERS_reg_16_33_inst : DFF_X1 port map( D => n3449, CK => n760, Q => 
                           REGISTERS_16_33_port, QN => n_2058);
   REGISTERS_reg_16_32_inst : DFF_X1 port map( D => n3448, CK => n761, Q => 
                           REGISTERS_16_32_port, QN => n_2059);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n3447, CK => n761, Q => 
                           REGISTERS_16_31_port, QN => n_2060);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n3446, CK => n761, Q => 
                           REGISTERS_16_30_port, QN => n_2061);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n3445, CK => n761, Q => 
                           REGISTERS_16_29_port, QN => n_2062);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n3444, CK => n761, Q => 
                           REGISTERS_16_28_port, QN => n_2063);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n3443, CK => n761, Q => 
                           REGISTERS_16_27_port, QN => n_2064);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n3442, CK => n761, Q => 
                           REGISTERS_16_26_port, QN => n_2065);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n3441, CK => n761, Q => 
                           REGISTERS_16_25_port, QN => n_2066);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n3440, CK => n761, Q => 
                           REGISTERS_16_24_port, QN => n_2067);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n3439, CK => n761, Q => 
                           REGISTERS_16_23_port, QN => n_2068);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n3438, CK => n761, Q => 
                           REGISTERS_16_22_port, QN => n_2069);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n3437, CK => n762, Q => 
                           REGISTERS_16_21_port, QN => n_2070);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n3436, CK => n762, Q => 
                           REGISTERS_16_20_port, QN => n_2071);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n3435, CK => n762, Q => 
                           REGISTERS_16_19_port, QN => n_2072);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n3434, CK => n762, Q => 
                           REGISTERS_16_18_port, QN => n_2073);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n3433, CK => n762, Q => 
                           REGISTERS_16_17_port, QN => n_2074);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n3432, CK => n762, Q => 
                           REGISTERS_16_16_port, QN => n_2075);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n3431, CK => n762, Q => 
                           REGISTERS_16_15_port, QN => n_2076);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n3430, CK => n762, Q => 
                           REGISTERS_16_14_port, QN => n_2077);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n3429, CK => n762, Q => 
                           REGISTERS_16_13_port, QN => n_2078);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n3428, CK => n762, Q => 
                           REGISTERS_16_12_port, QN => n_2079);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n3427, CK => n762, Q => 
                           REGISTERS_16_11_port, QN => n_2080);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n3426, CK => n763, Q => 
                           REGISTERS_16_10_port, QN => n_2081);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n3425, CK => n763, Q => 
                           REGISTERS_16_9_port, QN => n_2082);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n3424, CK => n763, Q => 
                           REGISTERS_16_8_port, QN => n_2083);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n3423, CK => n763, Q => 
                           REGISTERS_16_7_port, QN => n_2084);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n3422, CK => n763, Q => 
                           REGISTERS_16_6_port, QN => n_2085);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n3421, CK => n763, Q => 
                           REGISTERS_16_5_port, QN => n_2086);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n3420, CK => n763, Q => 
                           REGISTERS_16_4_port, QN => n_2087);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n3419, CK => n763, Q => 
                           REGISTERS_16_3_port, QN => n_2088);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n3418, CK => n763, Q => 
                           REGISTERS_16_2_port, QN => n_2089);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n3417, CK => n763, Q => 
                           REGISTERS_16_1_port, QN => n_2090);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n3416, CK => n763, Q => 
                           REGISTERS_16_0_port, QN => n_2091);
   REGISTERS_reg_17_63_inst : DFF_X1 port map( D => n3415, CK => n764, Q => 
                           REGISTERS_17_63_port, QN => n_2092);
   REGISTERS_reg_17_62_inst : DFF_X1 port map( D => n3414, CK => n764, Q => 
                           REGISTERS_17_62_port, QN => n_2093);
   REGISTERS_reg_17_61_inst : DFF_X1 port map( D => n3413, CK => n764, Q => 
                           REGISTERS_17_61_port, QN => n_2094);
   REGISTERS_reg_17_60_inst : DFF_X1 port map( D => n3412, CK => n764, Q => 
                           REGISTERS_17_60_port, QN => n_2095);
   REGISTERS_reg_17_59_inst : DFF_X1 port map( D => n3411, CK => n764, Q => 
                           REGISTERS_17_59_port, QN => n_2096);
   REGISTERS_reg_17_58_inst : DFF_X1 port map( D => n3410, CK => n764, Q => 
                           REGISTERS_17_58_port, QN => n_2097);
   REGISTERS_reg_17_57_inst : DFF_X1 port map( D => n3409, CK => n764, Q => 
                           REGISTERS_17_57_port, QN => n_2098);
   REGISTERS_reg_17_56_inst : DFF_X1 port map( D => n3408, CK => n764, Q => 
                           REGISTERS_17_56_port, QN => n_2099);
   REGISTERS_reg_17_55_inst : DFF_X1 port map( D => n3407, CK => n764, Q => 
                           REGISTERS_17_55_port, QN => n_2100);
   REGISTERS_reg_17_54_inst : DFF_X1 port map( D => n3406, CK => n764, Q => 
                           REGISTERS_17_54_port, QN => n_2101);
   REGISTERS_reg_17_53_inst : DFF_X1 port map( D => n3405, CK => n764, Q => 
                           REGISTERS_17_53_port, QN => n_2102);
   REGISTERS_reg_17_52_inst : DFF_X1 port map( D => n3404, CK => n765, Q => 
                           REGISTERS_17_52_port, QN => n_2103);
   REGISTERS_reg_17_51_inst : DFF_X1 port map( D => n3403, CK => n765, Q => 
                           REGISTERS_17_51_port, QN => n_2104);
   REGISTERS_reg_17_50_inst : DFF_X1 port map( D => n3402, CK => n765, Q => 
                           REGISTERS_17_50_port, QN => n_2105);
   REGISTERS_reg_17_49_inst : DFF_X1 port map( D => n3401, CK => n765, Q => 
                           REGISTERS_17_49_port, QN => n_2106);
   REGISTERS_reg_17_48_inst : DFF_X1 port map( D => n3400, CK => n765, Q => 
                           REGISTERS_17_48_port, QN => n_2107);
   REGISTERS_reg_17_47_inst : DFF_X1 port map( D => n3399, CK => n765, Q => 
                           REGISTERS_17_47_port, QN => n_2108);
   REGISTERS_reg_17_46_inst : DFF_X1 port map( D => n3398, CK => n765, Q => 
                           REGISTERS_17_46_port, QN => n_2109);
   REGISTERS_reg_17_45_inst : DFF_X1 port map( D => n3397, CK => n765, Q => 
                           REGISTERS_17_45_port, QN => n_2110);
   REGISTERS_reg_17_44_inst : DFF_X1 port map( D => n3396, CK => n765, Q => 
                           REGISTERS_17_44_port, QN => n_2111);
   REGISTERS_reg_17_43_inst : DFF_X1 port map( D => n3395, CK => n765, Q => 
                           REGISTERS_17_43_port, QN => n_2112);
   REGISTERS_reg_17_42_inst : DFF_X1 port map( D => n3394, CK => n765, Q => 
                           REGISTERS_17_42_port, QN => n_2113);
   REGISTERS_reg_17_41_inst : DFF_X1 port map( D => n3393, CK => n766, Q => 
                           REGISTERS_17_41_port, QN => n_2114);
   REGISTERS_reg_17_40_inst : DFF_X1 port map( D => n3392, CK => n766, Q => 
                           REGISTERS_17_40_port, QN => n_2115);
   REGISTERS_reg_17_39_inst : DFF_X1 port map( D => n3391, CK => n766, Q => 
                           REGISTERS_17_39_port, QN => n_2116);
   REGISTERS_reg_17_38_inst : DFF_X1 port map( D => n3390, CK => n766, Q => 
                           REGISTERS_17_38_port, QN => n_2117);
   REGISTERS_reg_17_37_inst : DFF_X1 port map( D => n3389, CK => n766, Q => 
                           REGISTERS_17_37_port, QN => n_2118);
   REGISTERS_reg_17_36_inst : DFF_X1 port map( D => n3388, CK => n766, Q => 
                           REGISTERS_17_36_port, QN => n_2119);
   REGISTERS_reg_17_35_inst : DFF_X1 port map( D => n3387, CK => n766, Q => 
                           REGISTERS_17_35_port, QN => n_2120);
   REGISTERS_reg_17_34_inst : DFF_X1 port map( D => n3386, CK => n766, Q => 
                           REGISTERS_17_34_port, QN => n_2121);
   REGISTERS_reg_17_33_inst : DFF_X1 port map( D => n3385, CK => n766, Q => 
                           REGISTERS_17_33_port, QN => n_2122);
   REGISTERS_reg_17_32_inst : DFF_X1 port map( D => n3384, CK => n766, Q => 
                           REGISTERS_17_32_port, QN => n_2123);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n3383, CK => n766, Q => 
                           REGISTERS_17_31_port, QN => n_2124);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n3382, CK => n767, Q => 
                           REGISTERS_17_30_port, QN => n_2125);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n3381, CK => n767, Q => 
                           REGISTERS_17_29_port, QN => n_2126);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n3380, CK => n767, Q => 
                           REGISTERS_17_28_port, QN => n_2127);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n3379, CK => n767, Q => 
                           REGISTERS_17_27_port, QN => n_2128);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n3378, CK => n767, Q => 
                           REGISTERS_17_26_port, QN => n_2129);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n3377, CK => n767, Q => 
                           REGISTERS_17_25_port, QN => n_2130);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n3376, CK => n767, Q => 
                           REGISTERS_17_24_port, QN => n_2131);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n3375, CK => n767, Q => 
                           REGISTERS_17_23_port, QN => n_2132);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n3374, CK => n767, Q => 
                           REGISTERS_17_22_port, QN => n_2133);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n3373, CK => n767, Q => 
                           REGISTERS_17_21_port, QN => n_2134);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n3372, CK => n767, Q => 
                           REGISTERS_17_20_port, QN => n_2135);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n3371, CK => n768, Q => 
                           REGISTERS_17_19_port, QN => n_2136);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n3370, CK => n768, Q => 
                           REGISTERS_17_18_port, QN => n_2137);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n3369, CK => n768, Q => 
                           REGISTERS_17_17_port, QN => n_2138);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n3368, CK => n768, Q => 
                           REGISTERS_17_16_port, QN => n_2139);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n3367, CK => n768, Q => 
                           REGISTERS_17_15_port, QN => n_2140);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n3366, CK => n768, Q => 
                           REGISTERS_17_14_port, QN => n_2141);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n3365, CK => n768, Q => 
                           REGISTERS_17_13_port, QN => n_2142);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n3364, CK => n768, Q => 
                           REGISTERS_17_12_port, QN => n_2143);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n3363, CK => n768, Q => 
                           REGISTERS_17_11_port, QN => n_2144);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n3362, CK => n768, Q => 
                           REGISTERS_17_10_port, QN => n_2145);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n3361, CK => n768, Q => 
                           REGISTERS_17_9_port, QN => n_2146);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n3360, CK => n769, Q => 
                           REGISTERS_17_8_port, QN => n_2147);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n3359, CK => n769, Q => 
                           REGISTERS_17_7_port, QN => n_2148);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n3358, CK => n769, Q => 
                           REGISTERS_17_6_port, QN => n_2149);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n3357, CK => n769, Q => 
                           REGISTERS_17_5_port, QN => n_2150);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n3356, CK => n769, Q => 
                           REGISTERS_17_4_port, QN => n_2151);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n3355, CK => n769, Q => 
                           REGISTERS_17_3_port, QN => n_2152);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n3354, CK => n769, Q => 
                           REGISTERS_17_2_port, QN => n_2153);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n3353, CK => n769, Q => 
                           REGISTERS_17_1_port, QN => n_2154);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n3352, CK => n769, Q => 
                           REGISTERS_17_0_port, QN => n_2155);
   REGISTERS_reg_18_63_inst : DFF_X1 port map( D => n3351, CK => n769, Q => 
                           REGISTERS_18_63_port, QN => n_2156);
   REGISTERS_reg_18_62_inst : DFF_X1 port map( D => n3350, CK => n769, Q => 
                           REGISTERS_18_62_port, QN => n_2157);
   REGISTERS_reg_18_61_inst : DFF_X1 port map( D => n3349, CK => n770, Q => 
                           REGISTERS_18_61_port, QN => n_2158);
   REGISTERS_reg_18_60_inst : DFF_X1 port map( D => n3348, CK => n770, Q => 
                           REGISTERS_18_60_port, QN => n_2159);
   REGISTERS_reg_18_59_inst : DFF_X1 port map( D => n3347, CK => n770, Q => 
                           REGISTERS_18_59_port, QN => n_2160);
   REGISTERS_reg_18_58_inst : DFF_X1 port map( D => n3346, CK => n770, Q => 
                           REGISTERS_18_58_port, QN => n_2161);
   REGISTERS_reg_18_57_inst : DFF_X1 port map( D => n3345, CK => n770, Q => 
                           REGISTERS_18_57_port, QN => n_2162);
   REGISTERS_reg_18_56_inst : DFF_X1 port map( D => n3344, CK => n770, Q => 
                           REGISTERS_18_56_port, QN => n_2163);
   REGISTERS_reg_18_55_inst : DFF_X1 port map( D => n3343, CK => n770, Q => 
                           REGISTERS_18_55_port, QN => n_2164);
   REGISTERS_reg_18_54_inst : DFF_X1 port map( D => n3342, CK => n770, Q => 
                           REGISTERS_18_54_port, QN => n_2165);
   REGISTERS_reg_18_53_inst : DFF_X1 port map( D => n3341, CK => n770, Q => 
                           REGISTERS_18_53_port, QN => n_2166);
   REGISTERS_reg_18_52_inst : DFF_X1 port map( D => n3340, CK => n770, Q => 
                           REGISTERS_18_52_port, QN => n_2167);
   REGISTERS_reg_18_51_inst : DFF_X1 port map( D => n3339, CK => n770, Q => 
                           REGISTERS_18_51_port, QN => n_2168);
   REGISTERS_reg_18_50_inst : DFF_X1 port map( D => n3338, CK => n771, Q => 
                           REGISTERS_18_50_port, QN => n_2169);
   REGISTERS_reg_18_49_inst : DFF_X1 port map( D => n3337, CK => n771, Q => 
                           REGISTERS_18_49_port, QN => n_2170);
   REGISTERS_reg_18_48_inst : DFF_X1 port map( D => n3336, CK => n771, Q => 
                           REGISTERS_18_48_port, QN => n_2171);
   REGISTERS_reg_18_47_inst : DFF_X1 port map( D => n3335, CK => n771, Q => 
                           REGISTERS_18_47_port, QN => n_2172);
   REGISTERS_reg_18_46_inst : DFF_X1 port map( D => n3334, CK => n771, Q => 
                           REGISTERS_18_46_port, QN => n_2173);
   REGISTERS_reg_18_45_inst : DFF_X1 port map( D => n3333, CK => n771, Q => 
                           REGISTERS_18_45_port, QN => n_2174);
   REGISTERS_reg_18_44_inst : DFF_X1 port map( D => n3332, CK => n771, Q => 
                           REGISTERS_18_44_port, QN => n_2175);
   REGISTERS_reg_18_43_inst : DFF_X1 port map( D => n3331, CK => n771, Q => 
                           REGISTERS_18_43_port, QN => n_2176);
   REGISTERS_reg_18_42_inst : DFF_X1 port map( D => n3330, CK => n771, Q => 
                           REGISTERS_18_42_port, QN => n_2177);
   REGISTERS_reg_18_41_inst : DFF_X1 port map( D => n3329, CK => n771, Q => 
                           REGISTERS_18_41_port, QN => n_2178);
   REGISTERS_reg_18_40_inst : DFF_X1 port map( D => n3328, CK => n771, Q => 
                           REGISTERS_18_40_port, QN => n_2179);
   REGISTERS_reg_18_39_inst : DFF_X1 port map( D => n3327, CK => n772, Q => 
                           REGISTERS_18_39_port, QN => n_2180);
   REGISTERS_reg_18_38_inst : DFF_X1 port map( D => n3326, CK => n772, Q => 
                           REGISTERS_18_38_port, QN => n_2181);
   REGISTERS_reg_18_37_inst : DFF_X1 port map( D => n3325, CK => n772, Q => 
                           REGISTERS_18_37_port, QN => n_2182);
   REGISTERS_reg_18_36_inst : DFF_X1 port map( D => n3324, CK => n772, Q => 
                           REGISTERS_18_36_port, QN => n_2183);
   REGISTERS_reg_18_35_inst : DFF_X1 port map( D => n3323, CK => n772, Q => 
                           REGISTERS_18_35_port, QN => n_2184);
   REGISTERS_reg_18_34_inst : DFF_X1 port map( D => n3322, CK => n772, Q => 
                           REGISTERS_18_34_port, QN => n_2185);
   REGISTERS_reg_18_33_inst : DFF_X1 port map( D => n3321, CK => n772, Q => 
                           REGISTERS_18_33_port, QN => n_2186);
   REGISTERS_reg_18_32_inst : DFF_X1 port map( D => n3320, CK => n772, Q => 
                           REGISTERS_18_32_port, QN => n_2187);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n3319, CK => n772, Q => 
                           REGISTERS_18_31_port, QN => n_2188);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n3318, CK => n772, Q => 
                           REGISTERS_18_30_port, QN => n_2189);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n3317, CK => n772, Q => 
                           REGISTERS_18_29_port, QN => n_2190);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n3316, CK => n773, Q => 
                           REGISTERS_18_28_port, QN => n_2191);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n3315, CK => n773, Q => 
                           REGISTERS_18_27_port, QN => n_2192);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n3314, CK => n773, Q => 
                           REGISTERS_18_26_port, QN => n_2193);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n3313, CK => n773, Q => 
                           REGISTERS_18_25_port, QN => n_2194);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n3312, CK => n773, Q => 
                           REGISTERS_18_24_port, QN => n_2195);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n3311, CK => n773, Q => 
                           REGISTERS_18_23_port, QN => n_2196);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n3310, CK => n773, Q => 
                           REGISTERS_18_22_port, QN => n_2197);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n3309, CK => n773, Q => 
                           REGISTERS_18_21_port, QN => n_2198);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n3308, CK => n773, Q => 
                           REGISTERS_18_20_port, QN => n_2199);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n3307, CK => n773, Q => 
                           REGISTERS_18_19_port, QN => n_2200);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n3306, CK => n773, Q => 
                           REGISTERS_18_18_port, QN => n_2201);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n3305, CK => n774, Q => 
                           REGISTERS_18_17_port, QN => n_2202);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n3304, CK => n774, Q => 
                           REGISTERS_18_16_port, QN => n_2203);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n3303, CK => n774, Q => 
                           REGISTERS_18_15_port, QN => n_2204);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n3302, CK => n774, Q => 
                           REGISTERS_18_14_port, QN => n_2205);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n3301, CK => n774, Q => 
                           REGISTERS_18_13_port, QN => n_2206);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n3300, CK => n774, Q => 
                           REGISTERS_18_12_port, QN => n_2207);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n3299, CK => n774, Q => 
                           REGISTERS_18_11_port, QN => n_2208);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n3298, CK => n774, Q => 
                           REGISTERS_18_10_port, QN => n_2209);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n3297, CK => n774, Q => 
                           REGISTERS_18_9_port, QN => n_2210);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n3296, CK => n774, Q => 
                           REGISTERS_18_8_port, QN => n_2211);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n3295, CK => n774, Q => 
                           REGISTERS_18_7_port, QN => n_2212);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n3294, CK => n775, Q => 
                           REGISTERS_18_6_port, QN => n_2213);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n3293, CK => n775, Q => 
                           REGISTERS_18_5_port, QN => n_2214);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n3292, CK => n775, Q => 
                           REGISTERS_18_4_port, QN => n_2215);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n3291, CK => n775, Q => 
                           REGISTERS_18_3_port, QN => n_2216);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n3290, CK => n775, Q => 
                           REGISTERS_18_2_port, QN => n_2217);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n3289, CK => n775, Q => 
                           REGISTERS_18_1_port, QN => n_2218);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n3288, CK => n775, Q => 
                           REGISTERS_18_0_port, QN => n_2219);
   REGISTERS_reg_19_63_inst : DFF_X1 port map( D => n3287, CK => n775, Q => 
                           REGISTERS_19_63_port, QN => n_2220);
   REGISTERS_reg_19_62_inst : DFF_X1 port map( D => n3286, CK => n775, Q => 
                           REGISTERS_19_62_port, QN => n_2221);
   REGISTERS_reg_19_61_inst : DFF_X1 port map( D => n3285, CK => n775, Q => 
                           REGISTERS_19_61_port, QN => n_2222);
   REGISTERS_reg_19_60_inst : DFF_X1 port map( D => n3284, CK => n775, Q => 
                           REGISTERS_19_60_port, QN => n_2223);
   REGISTERS_reg_19_59_inst : DFF_X1 port map( D => n3283, CK => n776, Q => 
                           REGISTERS_19_59_port, QN => n_2224);
   REGISTERS_reg_19_58_inst : DFF_X1 port map( D => n3282, CK => n776, Q => 
                           REGISTERS_19_58_port, QN => n_2225);
   REGISTERS_reg_19_57_inst : DFF_X1 port map( D => n3281, CK => n776, Q => 
                           REGISTERS_19_57_port, QN => n_2226);
   REGISTERS_reg_19_56_inst : DFF_X1 port map( D => n3280, CK => n776, Q => 
                           REGISTERS_19_56_port, QN => n_2227);
   REGISTERS_reg_19_55_inst : DFF_X1 port map( D => n3279, CK => n776, Q => 
                           REGISTERS_19_55_port, QN => n_2228);
   REGISTERS_reg_19_54_inst : DFF_X1 port map( D => n3278, CK => n776, Q => 
                           REGISTERS_19_54_port, QN => n_2229);
   REGISTERS_reg_19_53_inst : DFF_X1 port map( D => n3277, CK => n776, Q => 
                           REGISTERS_19_53_port, QN => n_2230);
   REGISTERS_reg_19_52_inst : DFF_X1 port map( D => n3276, CK => n776, Q => 
                           REGISTERS_19_52_port, QN => n_2231);
   REGISTERS_reg_19_51_inst : DFF_X1 port map( D => n3275, CK => n776, Q => 
                           REGISTERS_19_51_port, QN => n_2232);
   REGISTERS_reg_19_50_inst : DFF_X1 port map( D => n3274, CK => n776, Q => 
                           REGISTERS_19_50_port, QN => n_2233);
   REGISTERS_reg_19_49_inst : DFF_X1 port map( D => n3273, CK => n776, Q => 
                           REGISTERS_19_49_port, QN => n_2234);
   REGISTERS_reg_19_48_inst : DFF_X1 port map( D => n3272, CK => n777, Q => 
                           REGISTERS_19_48_port, QN => n_2235);
   REGISTERS_reg_19_47_inst : DFF_X1 port map( D => n3271, CK => n777, Q => 
                           REGISTERS_19_47_port, QN => n_2236);
   REGISTERS_reg_19_46_inst : DFF_X1 port map( D => n3270, CK => n777, Q => 
                           REGISTERS_19_46_port, QN => n_2237);
   REGISTERS_reg_19_45_inst : DFF_X1 port map( D => n3269, CK => n777, Q => 
                           REGISTERS_19_45_port, QN => n_2238);
   REGISTERS_reg_19_44_inst : DFF_X1 port map( D => n3268, CK => n777, Q => 
                           REGISTERS_19_44_port, QN => n_2239);
   REGISTERS_reg_19_43_inst : DFF_X1 port map( D => n3267, CK => n777, Q => 
                           REGISTERS_19_43_port, QN => n_2240);
   REGISTERS_reg_19_42_inst : DFF_X1 port map( D => n3266, CK => n777, Q => 
                           REGISTERS_19_42_port, QN => n_2241);
   REGISTERS_reg_19_41_inst : DFF_X1 port map( D => n3265, CK => n777, Q => 
                           REGISTERS_19_41_port, QN => n_2242);
   REGISTERS_reg_19_40_inst : DFF_X1 port map( D => n3264, CK => n777, Q => 
                           REGISTERS_19_40_port, QN => n_2243);
   REGISTERS_reg_19_39_inst : DFF_X1 port map( D => n3263, CK => n777, Q => 
                           REGISTERS_19_39_port, QN => n_2244);
   REGISTERS_reg_19_38_inst : DFF_X1 port map( D => n3262, CK => n777, Q => 
                           REGISTERS_19_38_port, QN => n_2245);
   REGISTERS_reg_19_37_inst : DFF_X1 port map( D => n3261, CK => n778, Q => 
                           REGISTERS_19_37_port, QN => n_2246);
   REGISTERS_reg_19_36_inst : DFF_X1 port map( D => n3260, CK => n778, Q => 
                           REGISTERS_19_36_port, QN => n_2247);
   REGISTERS_reg_19_35_inst : DFF_X1 port map( D => n3259, CK => n778, Q => 
                           REGISTERS_19_35_port, QN => n_2248);
   REGISTERS_reg_19_34_inst : DFF_X1 port map( D => n3258, CK => n778, Q => 
                           REGISTERS_19_34_port, QN => n_2249);
   REGISTERS_reg_19_33_inst : DFF_X1 port map( D => n3257, CK => n778, Q => 
                           REGISTERS_19_33_port, QN => n_2250);
   REGISTERS_reg_19_32_inst : DFF_X1 port map( D => n3256, CK => n778, Q => 
                           REGISTERS_19_32_port, QN => n_2251);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n3255, CK => n778, Q => 
                           REGISTERS_19_31_port, QN => n_2252);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n3254, CK => n778, Q => 
                           REGISTERS_19_30_port, QN => n_2253);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n3253, CK => n778, Q => 
                           REGISTERS_19_29_port, QN => n_2254);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n3252, CK => n778, Q => 
                           REGISTERS_19_28_port, QN => n_2255);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n3251, CK => n778, Q => 
                           REGISTERS_19_27_port, QN => n_2256);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n3250, CK => n779, Q => 
                           REGISTERS_19_26_port, QN => n_2257);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n3249, CK => n779, Q => 
                           REGISTERS_19_25_port, QN => n_2258);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n3248, CK => n779, Q => 
                           REGISTERS_19_24_port, QN => n_2259);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n3247, CK => n779, Q => 
                           REGISTERS_19_23_port, QN => n_2260);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n3246, CK => n779, Q => 
                           REGISTERS_19_22_port, QN => n_2261);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n3245, CK => n779, Q => 
                           REGISTERS_19_21_port, QN => n_2262);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n3244, CK => n779, Q => 
                           REGISTERS_19_20_port, QN => n_2263);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n3243, CK => n779, Q => 
                           REGISTERS_19_19_port, QN => n_2264);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n3242, CK => n779, Q => 
                           REGISTERS_19_18_port, QN => n_2265);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n3241, CK => n779, Q => 
                           REGISTERS_19_17_port, QN => n_2266);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n3240, CK => n779, Q => 
                           REGISTERS_19_16_port, QN => n_2267);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n3239, CK => n780, Q => 
                           REGISTERS_19_15_port, QN => n_2268);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n3238, CK => n780, Q => 
                           REGISTERS_19_14_port, QN => n_2269);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n3237, CK => n780, Q => 
                           REGISTERS_19_13_port, QN => n_2270);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n3236, CK => n780, Q => 
                           REGISTERS_19_12_port, QN => n_2271);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n3235, CK => n780, Q => 
                           REGISTERS_19_11_port, QN => n_2272);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n3234, CK => n780, Q => 
                           REGISTERS_19_10_port, QN => n_2273);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n3233, CK => n780, Q => 
                           REGISTERS_19_9_port, QN => n_2274);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n3232, CK => n780, Q => 
                           REGISTERS_19_8_port, QN => n_2275);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n3231, CK => n780, Q => 
                           REGISTERS_19_7_port, QN => n_2276);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n3230, CK => n780, Q => 
                           REGISTERS_19_6_port, QN => n_2277);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n3229, CK => n780, Q => 
                           REGISTERS_19_5_port, QN => n_2278);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n3228, CK => n781, Q => 
                           REGISTERS_19_4_port, QN => n_2279);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n3227, CK => n781, Q => 
                           REGISTERS_19_3_port, QN => n_2280);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n3226, CK => n781, Q => 
                           REGISTERS_19_2_port, QN => n_2281);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n3225, CK => n781, Q => 
                           REGISTERS_19_1_port, QN => n_2282);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n3224, CK => n781, Q => 
                           REGISTERS_19_0_port, QN => n_2283);
   REGISTERS_reg_20_63_inst : DFF_X1 port map( D => n3223, CK => n781, Q => 
                           REGISTERS_20_63_port, QN => n_2284);
   REGISTERS_reg_20_62_inst : DFF_X1 port map( D => n3222, CK => n781, Q => 
                           REGISTERS_20_62_port, QN => n_2285);
   REGISTERS_reg_20_61_inst : DFF_X1 port map( D => n3221, CK => n781, Q => 
                           REGISTERS_20_61_port, QN => n_2286);
   REGISTERS_reg_20_60_inst : DFF_X1 port map( D => n3220, CK => n781, Q => 
                           REGISTERS_20_60_port, QN => n_2287);
   REGISTERS_reg_20_59_inst : DFF_X1 port map( D => n3219, CK => n781, Q => 
                           REGISTERS_20_59_port, QN => n_2288);
   REGISTERS_reg_20_58_inst : DFF_X1 port map( D => n3218, CK => n781, Q => 
                           REGISTERS_20_58_port, QN => n_2289);
   REGISTERS_reg_20_57_inst : DFF_X1 port map( D => n3217, CK => n782, Q => 
                           REGISTERS_20_57_port, QN => n_2290);
   REGISTERS_reg_20_56_inst : DFF_X1 port map( D => n3216, CK => n782, Q => 
                           REGISTERS_20_56_port, QN => n_2291);
   REGISTERS_reg_20_55_inst : DFF_X1 port map( D => n3215, CK => n782, Q => 
                           REGISTERS_20_55_port, QN => n_2292);
   REGISTERS_reg_20_54_inst : DFF_X1 port map( D => n3214, CK => n782, Q => 
                           REGISTERS_20_54_port, QN => n_2293);
   REGISTERS_reg_20_53_inst : DFF_X1 port map( D => n3213, CK => n782, Q => 
                           REGISTERS_20_53_port, QN => n_2294);
   REGISTERS_reg_20_52_inst : DFF_X1 port map( D => n3212, CK => n782, Q => 
                           REGISTERS_20_52_port, QN => n_2295);
   REGISTERS_reg_20_51_inst : DFF_X1 port map( D => n3211, CK => n782, Q => 
                           REGISTERS_20_51_port, QN => n_2296);
   REGISTERS_reg_20_50_inst : DFF_X1 port map( D => n3210, CK => n782, Q => 
                           REGISTERS_20_50_port, QN => n_2297);
   REGISTERS_reg_20_49_inst : DFF_X1 port map( D => n3209, CK => n782, Q => 
                           REGISTERS_20_49_port, QN => n_2298);
   REGISTERS_reg_20_48_inst : DFF_X1 port map( D => n3208, CK => n782, Q => 
                           REGISTERS_20_48_port, QN => n_2299);
   REGISTERS_reg_20_47_inst : DFF_X1 port map( D => n3207, CK => n782, Q => 
                           REGISTERS_20_47_port, QN => n_2300);
   REGISTERS_reg_20_46_inst : DFF_X1 port map( D => n3206, CK => n783, Q => 
                           REGISTERS_20_46_port, QN => n_2301);
   REGISTERS_reg_20_45_inst : DFF_X1 port map( D => n3205, CK => n783, Q => 
                           REGISTERS_20_45_port, QN => n_2302);
   REGISTERS_reg_20_44_inst : DFF_X1 port map( D => n3204, CK => n783, Q => 
                           REGISTERS_20_44_port, QN => n_2303);
   REGISTERS_reg_20_43_inst : DFF_X1 port map( D => n3203, CK => n783, Q => 
                           REGISTERS_20_43_port, QN => n_2304);
   REGISTERS_reg_20_42_inst : DFF_X1 port map( D => n3202, CK => n783, Q => 
                           REGISTERS_20_42_port, QN => n_2305);
   REGISTERS_reg_20_41_inst : DFF_X1 port map( D => n3201, CK => n783, Q => 
                           REGISTERS_20_41_port, QN => n_2306);
   REGISTERS_reg_20_40_inst : DFF_X1 port map( D => n3200, CK => n783, Q => 
                           REGISTERS_20_40_port, QN => n_2307);
   REGISTERS_reg_20_39_inst : DFF_X1 port map( D => n3199, CK => n783, Q => 
                           REGISTERS_20_39_port, QN => n_2308);
   REGISTERS_reg_20_38_inst : DFF_X1 port map( D => n3198, CK => n783, Q => 
                           REGISTERS_20_38_port, QN => n_2309);
   REGISTERS_reg_20_37_inst : DFF_X1 port map( D => n3197, CK => n783, Q => 
                           REGISTERS_20_37_port, QN => n_2310);
   REGISTERS_reg_20_36_inst : DFF_X1 port map( D => n3196, CK => n783, Q => 
                           REGISTERS_20_36_port, QN => n_2311);
   REGISTERS_reg_20_35_inst : DFF_X1 port map( D => n3195, CK => n784, Q => 
                           REGISTERS_20_35_port, QN => n_2312);
   REGISTERS_reg_20_34_inst : DFF_X1 port map( D => n3194, CK => n784, Q => 
                           REGISTERS_20_34_port, QN => n_2313);
   REGISTERS_reg_20_33_inst : DFF_X1 port map( D => n3193, CK => n784, Q => 
                           REGISTERS_20_33_port, QN => n_2314);
   REGISTERS_reg_20_32_inst : DFF_X1 port map( D => n3192, CK => n784, Q => 
                           REGISTERS_20_32_port, QN => n_2315);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n3191, CK => n784, Q => 
                           REGISTERS_20_31_port, QN => n_2316);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n3190, CK => n784, Q => 
                           REGISTERS_20_30_port, QN => n_2317);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n3189, CK => n784, Q => 
                           REGISTERS_20_29_port, QN => n_2318);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n3188, CK => n784, Q => 
                           REGISTERS_20_28_port, QN => n_2319);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n3187, CK => n784, Q => 
                           REGISTERS_20_27_port, QN => n_2320);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n3186, CK => n784, Q => 
                           REGISTERS_20_26_port, QN => n_2321);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n3185, CK => n784, Q => 
                           REGISTERS_20_25_port, QN => n_2322);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n3184, CK => n785, Q => 
                           REGISTERS_20_24_port, QN => n_2323);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n3183, CK => n785, Q => 
                           REGISTERS_20_23_port, QN => n_2324);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n3182, CK => n785, Q => 
                           REGISTERS_20_22_port, QN => n_2325);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n3181, CK => n785, Q => 
                           REGISTERS_20_21_port, QN => n_2326);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n3180, CK => n785, Q => 
                           REGISTERS_20_20_port, QN => n_2327);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n3179, CK => n785, Q => 
                           REGISTERS_20_19_port, QN => n_2328);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n3178, CK => n785, Q => 
                           REGISTERS_20_18_port, QN => n_2329);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n3177, CK => n785, Q => 
                           REGISTERS_20_17_port, QN => n_2330);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n3176, CK => n785, Q => 
                           REGISTERS_20_16_port, QN => n_2331);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n3175, CK => n785, Q => 
                           REGISTERS_20_15_port, QN => n_2332);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n3174, CK => n785, Q => 
                           REGISTERS_20_14_port, QN => n_2333);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n3173, CK => n786, Q => 
                           REGISTERS_20_13_port, QN => n_2334);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n3172, CK => n786, Q => 
                           REGISTERS_20_12_port, QN => n_2335);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n3171, CK => n786, Q => 
                           REGISTERS_20_11_port, QN => n_2336);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n3170, CK => n786, Q => 
                           REGISTERS_20_10_port, QN => n_2337);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n3169, CK => n786, Q => 
                           REGISTERS_20_9_port, QN => n_2338);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n3168, CK => n786, Q => 
                           REGISTERS_20_8_port, QN => n_2339);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n3167, CK => n786, Q => 
                           REGISTERS_20_7_port, QN => n_2340);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n3166, CK => n786, Q => 
                           REGISTERS_20_6_port, QN => n_2341);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n3165, CK => n786, Q => 
                           REGISTERS_20_5_port, QN => n_2342);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n3164, CK => n786, Q => 
                           REGISTERS_20_4_port, QN => n_2343);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n3163, CK => n786, Q => 
                           REGISTERS_20_3_port, QN => n_2344);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n3162, CK => n787, Q => 
                           REGISTERS_20_2_port, QN => n_2345);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n3161, CK => n787, Q => 
                           REGISTERS_20_1_port, QN => n_2346);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n3160, CK => n787, Q => 
                           REGISTERS_20_0_port, QN => n_2347);
   REGISTERS_reg_21_63_inst : DFF_X1 port map( D => n3159, CK => n787, Q => 
                           REGISTERS_21_63_port, QN => n_2348);
   REGISTERS_reg_21_62_inst : DFF_X1 port map( D => n3158, CK => n787, Q => 
                           REGISTERS_21_62_port, QN => n_2349);
   REGISTERS_reg_21_61_inst : DFF_X1 port map( D => n3157, CK => n787, Q => 
                           REGISTERS_21_61_port, QN => n_2350);
   REGISTERS_reg_21_60_inst : DFF_X1 port map( D => n3156, CK => n787, Q => 
                           REGISTERS_21_60_port, QN => n_2351);
   REGISTERS_reg_21_59_inst : DFF_X1 port map( D => n3155, CK => n787, Q => 
                           REGISTERS_21_59_port, QN => n_2352);
   REGISTERS_reg_21_58_inst : DFF_X1 port map( D => n3154, CK => n787, Q => 
                           REGISTERS_21_58_port, QN => n_2353);
   REGISTERS_reg_21_57_inst : DFF_X1 port map( D => n3153, CK => n787, Q => 
                           REGISTERS_21_57_port, QN => n_2354);
   REGISTERS_reg_21_56_inst : DFF_X1 port map( D => n3152, CK => n787, Q => 
                           REGISTERS_21_56_port, QN => n_2355);
   REGISTERS_reg_21_55_inst : DFF_X1 port map( D => n3151, CK => n788, Q => 
                           REGISTERS_21_55_port, QN => n_2356);
   REGISTERS_reg_21_54_inst : DFF_X1 port map( D => n3150, CK => n788, Q => 
                           REGISTERS_21_54_port, QN => n_2357);
   REGISTERS_reg_21_53_inst : DFF_X1 port map( D => n3149, CK => n788, Q => 
                           REGISTERS_21_53_port, QN => n_2358);
   REGISTERS_reg_21_52_inst : DFF_X1 port map( D => n3148, CK => n788, Q => 
                           REGISTERS_21_52_port, QN => n_2359);
   REGISTERS_reg_21_51_inst : DFF_X1 port map( D => n3147, CK => n788, Q => 
                           REGISTERS_21_51_port, QN => n_2360);
   REGISTERS_reg_21_50_inst : DFF_X1 port map( D => n3146, CK => n788, Q => 
                           REGISTERS_21_50_port, QN => n_2361);
   REGISTERS_reg_21_49_inst : DFF_X1 port map( D => n3145, CK => n788, Q => 
                           REGISTERS_21_49_port, QN => n_2362);
   REGISTERS_reg_21_48_inst : DFF_X1 port map( D => n3144, CK => n788, Q => 
                           REGISTERS_21_48_port, QN => n_2363);
   REGISTERS_reg_21_47_inst : DFF_X1 port map( D => n3143, CK => n788, Q => 
                           REGISTERS_21_47_port, QN => n_2364);
   REGISTERS_reg_21_46_inst : DFF_X1 port map( D => n3142, CK => n788, Q => 
                           REGISTERS_21_46_port, QN => n_2365);
   REGISTERS_reg_21_45_inst : DFF_X1 port map( D => n3141, CK => n788, Q => 
                           REGISTERS_21_45_port, QN => n_2366);
   REGISTERS_reg_21_44_inst : DFF_X1 port map( D => n3140, CK => n789, Q => 
                           REGISTERS_21_44_port, QN => n_2367);
   REGISTERS_reg_21_43_inst : DFF_X1 port map( D => n3139, CK => n789, Q => 
                           REGISTERS_21_43_port, QN => n_2368);
   REGISTERS_reg_21_42_inst : DFF_X1 port map( D => n3138, CK => n789, Q => 
                           REGISTERS_21_42_port, QN => n_2369);
   REGISTERS_reg_21_41_inst : DFF_X1 port map( D => n3137, CK => n789, Q => 
                           REGISTERS_21_41_port, QN => n_2370);
   REGISTERS_reg_21_40_inst : DFF_X1 port map( D => n3136, CK => n789, Q => 
                           REGISTERS_21_40_port, QN => n_2371);
   REGISTERS_reg_21_39_inst : DFF_X1 port map( D => n3135, CK => n789, Q => 
                           REGISTERS_21_39_port, QN => n_2372);
   REGISTERS_reg_21_38_inst : DFF_X1 port map( D => n3134, CK => n789, Q => 
                           REGISTERS_21_38_port, QN => n_2373);
   REGISTERS_reg_21_37_inst : DFF_X1 port map( D => n3133, CK => n789, Q => 
                           REGISTERS_21_37_port, QN => n_2374);
   REGISTERS_reg_21_36_inst : DFF_X1 port map( D => n3132, CK => n789, Q => 
                           REGISTERS_21_36_port, QN => n_2375);
   REGISTERS_reg_21_35_inst : DFF_X1 port map( D => n3131, CK => n789, Q => 
                           REGISTERS_21_35_port, QN => n_2376);
   REGISTERS_reg_21_34_inst : DFF_X1 port map( D => n3130, CK => n789, Q => 
                           REGISTERS_21_34_port, QN => n_2377);
   REGISTERS_reg_21_33_inst : DFF_X1 port map( D => n3129, CK => n790, Q => 
                           REGISTERS_21_33_port, QN => n_2378);
   REGISTERS_reg_21_32_inst : DFF_X1 port map( D => n3128, CK => n790, Q => 
                           REGISTERS_21_32_port, QN => n_2379);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n3127, CK => n790, Q => 
                           REGISTERS_21_31_port, QN => n_2380);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n3126, CK => n790, Q => 
                           REGISTERS_21_30_port, QN => n_2381);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n3125, CK => n790, Q => 
                           REGISTERS_21_29_port, QN => n_2382);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n3124, CK => n790, Q => 
                           REGISTERS_21_28_port, QN => n_2383);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n3123, CK => n790, Q => 
                           REGISTERS_21_27_port, QN => n_2384);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n3122, CK => n790, Q => 
                           REGISTERS_21_26_port, QN => n_2385);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n3121, CK => n790, Q => 
                           REGISTERS_21_25_port, QN => n_2386);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n3120, CK => n790, Q => 
                           REGISTERS_21_24_port, QN => n_2387);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n3119, CK => n790, Q => 
                           REGISTERS_21_23_port, QN => n_2388);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n3118, CK => n791, Q => 
                           REGISTERS_21_22_port, QN => n_2389);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n3117, CK => n791, Q => 
                           REGISTERS_21_21_port, QN => n_2390);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n3116, CK => n791, Q => 
                           REGISTERS_21_20_port, QN => n_2391);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n3115, CK => n791, Q => 
                           REGISTERS_21_19_port, QN => n_2392);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n3114, CK => n791, Q => 
                           REGISTERS_21_18_port, QN => n_2393);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n3113, CK => n791, Q => 
                           REGISTERS_21_17_port, QN => n_2394);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n3112, CK => n791, Q => 
                           REGISTERS_21_16_port, QN => n_2395);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n3111, CK => n791, Q => 
                           REGISTERS_21_15_port, QN => n_2396);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n3110, CK => n791, Q => 
                           REGISTERS_21_14_port, QN => n_2397);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n3109, CK => n791, Q => 
                           REGISTERS_21_13_port, QN => n_2398);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n3108, CK => n791, Q => 
                           REGISTERS_21_12_port, QN => n_2399);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n3107, CK => n792, Q => 
                           REGISTERS_21_11_port, QN => n_2400);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n3106, CK => n792, Q => 
                           REGISTERS_21_10_port, QN => n_2401);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n3105, CK => n792, Q => 
                           REGISTERS_21_9_port, QN => n_2402);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n3104, CK => n792, Q => 
                           REGISTERS_21_8_port, QN => n_2403);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n3103, CK => n792, Q => 
                           REGISTERS_21_7_port, QN => n_2404);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n3102, CK => n792, Q => 
                           REGISTERS_21_6_port, QN => n_2405);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n3101, CK => n792, Q => 
                           REGISTERS_21_5_port, QN => n_2406);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n3100, CK => n792, Q => 
                           REGISTERS_21_4_port, QN => n_2407);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n3099, CK => n792, Q => 
                           REGISTERS_21_3_port, QN => n_2408);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n3098, CK => n792, Q => 
                           REGISTERS_21_2_port, QN => n_2409);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n3097, CK => n792, Q => 
                           REGISTERS_21_1_port, QN => n_2410);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n3096, CK => n793, Q => 
                           REGISTERS_21_0_port, QN => n_2411);
   REGISTERS_reg_22_63_inst : DFF_X1 port map( D => n3095, CK => n793, Q => 
                           REGISTERS_22_63_port, QN => n_2412);
   REGISTERS_reg_22_62_inst : DFF_X1 port map( D => n3094, CK => n793, Q => 
                           REGISTERS_22_62_port, QN => n_2413);
   REGISTERS_reg_22_61_inst : DFF_X1 port map( D => n3093, CK => n793, Q => 
                           REGISTERS_22_61_port, QN => n_2414);
   REGISTERS_reg_22_60_inst : DFF_X1 port map( D => n3092, CK => n793, Q => 
                           REGISTERS_22_60_port, QN => n_2415);
   REGISTERS_reg_22_59_inst : DFF_X1 port map( D => n3091, CK => n793, Q => 
                           REGISTERS_22_59_port, QN => n_2416);
   REGISTERS_reg_22_58_inst : DFF_X1 port map( D => n3090, CK => n793, Q => 
                           REGISTERS_22_58_port, QN => n_2417);
   REGISTERS_reg_22_57_inst : DFF_X1 port map( D => n3089, CK => n793, Q => 
                           REGISTERS_22_57_port, QN => n_2418);
   REGISTERS_reg_22_56_inst : DFF_X1 port map( D => n3088, CK => n793, Q => 
                           REGISTERS_22_56_port, QN => n_2419);
   REGISTERS_reg_22_55_inst : DFF_X1 port map( D => n3087, CK => n793, Q => 
                           REGISTERS_22_55_port, QN => n_2420);
   REGISTERS_reg_22_54_inst : DFF_X1 port map( D => n3086, CK => n793, Q => 
                           REGISTERS_22_54_port, QN => n_2421);
   REGISTERS_reg_22_53_inst : DFF_X1 port map( D => n3085, CK => n794, Q => 
                           REGISTERS_22_53_port, QN => n_2422);
   REGISTERS_reg_22_52_inst : DFF_X1 port map( D => n3084, CK => n794, Q => 
                           REGISTERS_22_52_port, QN => n_2423);
   REGISTERS_reg_22_51_inst : DFF_X1 port map( D => n3083, CK => n794, Q => 
                           REGISTERS_22_51_port, QN => n_2424);
   REGISTERS_reg_22_50_inst : DFF_X1 port map( D => n3082, CK => n794, Q => 
                           REGISTERS_22_50_port, QN => n_2425);
   REGISTERS_reg_22_49_inst : DFF_X1 port map( D => n3081, CK => n794, Q => 
                           REGISTERS_22_49_port, QN => n_2426);
   REGISTERS_reg_22_48_inst : DFF_X1 port map( D => n3080, CK => n794, Q => 
                           REGISTERS_22_48_port, QN => n_2427);
   REGISTERS_reg_22_47_inst : DFF_X1 port map( D => n3079, CK => n794, Q => 
                           REGISTERS_22_47_port, QN => n_2428);
   REGISTERS_reg_22_46_inst : DFF_X1 port map( D => n3078, CK => n794, Q => 
                           REGISTERS_22_46_port, QN => n_2429);
   REGISTERS_reg_22_45_inst : DFF_X1 port map( D => n3077, CK => n794, Q => 
                           REGISTERS_22_45_port, QN => n_2430);
   REGISTERS_reg_22_44_inst : DFF_X1 port map( D => n3076, CK => n794, Q => 
                           REGISTERS_22_44_port, QN => n_2431);
   REGISTERS_reg_22_43_inst : DFF_X1 port map( D => n3075, CK => n794, Q => 
                           REGISTERS_22_43_port, QN => n_2432);
   REGISTERS_reg_22_42_inst : DFF_X1 port map( D => n3074, CK => n795, Q => 
                           REGISTERS_22_42_port, QN => n_2433);
   REGISTERS_reg_22_41_inst : DFF_X1 port map( D => n3073, CK => n795, Q => 
                           REGISTERS_22_41_port, QN => n_2434);
   REGISTERS_reg_22_40_inst : DFF_X1 port map( D => n3072, CK => n795, Q => 
                           REGISTERS_22_40_port, QN => n_2435);
   REGISTERS_reg_22_39_inst : DFF_X1 port map( D => n3071, CK => n795, Q => 
                           REGISTERS_22_39_port, QN => n_2436);
   REGISTERS_reg_22_38_inst : DFF_X1 port map( D => n3070, CK => n795, Q => 
                           REGISTERS_22_38_port, QN => n_2437);
   REGISTERS_reg_22_37_inst : DFF_X1 port map( D => n3069, CK => n795, Q => 
                           REGISTERS_22_37_port, QN => n_2438);
   REGISTERS_reg_22_36_inst : DFF_X1 port map( D => n3068, CK => n795, Q => 
                           REGISTERS_22_36_port, QN => n_2439);
   REGISTERS_reg_22_35_inst : DFF_X1 port map( D => n3067, CK => n795, Q => 
                           REGISTERS_22_35_port, QN => n_2440);
   REGISTERS_reg_22_34_inst : DFF_X1 port map( D => n3066, CK => n795, Q => 
                           REGISTERS_22_34_port, QN => n_2441);
   REGISTERS_reg_22_33_inst : DFF_X1 port map( D => n3065, CK => n795, Q => 
                           REGISTERS_22_33_port, QN => n_2442);
   REGISTERS_reg_22_32_inst : DFF_X1 port map( D => n3064, CK => n795, Q => 
                           REGISTERS_22_32_port, QN => n_2443);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n3063, CK => n796, Q => 
                           REGISTERS_22_31_port, QN => n_2444);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n3062, CK => n796, Q => 
                           REGISTERS_22_30_port, QN => n_2445);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n3061, CK => n796, Q => 
                           REGISTERS_22_29_port, QN => n_2446);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n3060, CK => n796, Q => 
                           REGISTERS_22_28_port, QN => n_2447);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n3059, CK => n796, Q => 
                           REGISTERS_22_27_port, QN => n_2448);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n3058, CK => n796, Q => 
                           REGISTERS_22_26_port, QN => n_2449);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n3057, CK => n796, Q => 
                           REGISTERS_22_25_port, QN => n_2450);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n3056, CK => n796, Q => 
                           REGISTERS_22_24_port, QN => n_2451);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n3055, CK => n796, Q => 
                           REGISTERS_22_23_port, QN => n_2452);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n3054, CK => n796, Q => 
                           REGISTERS_22_22_port, QN => n_2453);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n3053, CK => n796, Q => 
                           REGISTERS_22_21_port, QN => n_2454);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n3052, CK => n797, Q => 
                           REGISTERS_22_20_port, QN => n_2455);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n3051, CK => n797, Q => 
                           REGISTERS_22_19_port, QN => n_2456);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n3050, CK => n797, Q => 
                           REGISTERS_22_18_port, QN => n_2457);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n3049, CK => n797, Q => 
                           REGISTERS_22_17_port, QN => n_2458);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n3048, CK => n797, Q => 
                           REGISTERS_22_16_port, QN => n_2459);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n3047, CK => n797, Q => 
                           REGISTERS_22_15_port, QN => n_2460);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n3046, CK => n797, Q => 
                           REGISTERS_22_14_port, QN => n_2461);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n3045, CK => n797, Q => 
                           REGISTERS_22_13_port, QN => n_2462);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n3044, CK => n797, Q => 
                           REGISTERS_22_12_port, QN => n_2463);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n3043, CK => n797, Q => 
                           REGISTERS_22_11_port, QN => n_2464);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n3042, CK => n797, Q => 
                           REGISTERS_22_10_port, QN => n_2465);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n3041, CK => n798, Q => 
                           REGISTERS_22_9_port, QN => n_2466);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n3040, CK => n798, Q => 
                           REGISTERS_22_8_port, QN => n_2467);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n3039, CK => n798, Q => 
                           REGISTERS_22_7_port, QN => n_2468);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n3038, CK => n798, Q => 
                           REGISTERS_22_6_port, QN => n_2469);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n3037, CK => n798, Q => 
                           REGISTERS_22_5_port, QN => n_2470);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n3036, CK => n798, Q => 
                           REGISTERS_22_4_port, QN => n_2471);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n3035, CK => n798, Q => 
                           REGISTERS_22_3_port, QN => n_2472);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n3034, CK => n798, Q => 
                           REGISTERS_22_2_port, QN => n_2473);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n3033, CK => n798, Q => 
                           REGISTERS_22_1_port, QN => n_2474);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n3032, CK => n798, Q => 
                           REGISTERS_22_0_port, QN => n_2475);
   REGISTERS_reg_23_63_inst : DFF_X1 port map( D => n3031, CK => n798, Q => 
                           REGISTERS_23_63_port, QN => n_2476);
   REGISTERS_reg_23_62_inst : DFF_X1 port map( D => n3030, CK => n799, Q => 
                           REGISTERS_23_62_port, QN => n_2477);
   REGISTERS_reg_23_61_inst : DFF_X1 port map( D => n3029, CK => n799, Q => 
                           REGISTERS_23_61_port, QN => n_2478);
   REGISTERS_reg_23_60_inst : DFF_X1 port map( D => n3028, CK => n799, Q => 
                           REGISTERS_23_60_port, QN => n_2479);
   REGISTERS_reg_23_59_inst : DFF_X1 port map( D => n3027, CK => n799, Q => 
                           REGISTERS_23_59_port, QN => n_2480);
   REGISTERS_reg_23_58_inst : DFF_X1 port map( D => n3026, CK => n799, Q => 
                           REGISTERS_23_58_port, QN => n_2481);
   REGISTERS_reg_23_57_inst : DFF_X1 port map( D => n3025, CK => n799, Q => 
                           REGISTERS_23_57_port, QN => n_2482);
   REGISTERS_reg_23_56_inst : DFF_X1 port map( D => n3024, CK => n799, Q => 
                           REGISTERS_23_56_port, QN => n_2483);
   REGISTERS_reg_23_55_inst : DFF_X1 port map( D => n3023, CK => n799, Q => 
                           REGISTERS_23_55_port, QN => n_2484);
   REGISTERS_reg_23_54_inst : DFF_X1 port map( D => n3022, CK => n799, Q => 
                           REGISTERS_23_54_port, QN => n_2485);
   REGISTERS_reg_23_53_inst : DFF_X1 port map( D => n3021, CK => n799, Q => 
                           REGISTERS_23_53_port, QN => n_2486);
   REGISTERS_reg_23_52_inst : DFF_X1 port map( D => n3020, CK => n799, Q => 
                           REGISTERS_23_52_port, QN => n_2487);
   REGISTERS_reg_23_51_inst : DFF_X1 port map( D => n3019, CK => n800, Q => 
                           REGISTERS_23_51_port, QN => n_2488);
   REGISTERS_reg_23_50_inst : DFF_X1 port map( D => n3018, CK => n800, Q => 
                           REGISTERS_23_50_port, QN => n_2489);
   REGISTERS_reg_23_49_inst : DFF_X1 port map( D => n3017, CK => n800, Q => 
                           REGISTERS_23_49_port, QN => n_2490);
   REGISTERS_reg_23_48_inst : DFF_X1 port map( D => n3016, CK => n800, Q => 
                           REGISTERS_23_48_port, QN => n_2491);
   REGISTERS_reg_23_47_inst : DFF_X1 port map( D => n3015, CK => n800, Q => 
                           REGISTERS_23_47_port, QN => n_2492);
   REGISTERS_reg_23_46_inst : DFF_X1 port map( D => n3014, CK => n800, Q => 
                           REGISTERS_23_46_port, QN => n_2493);
   REGISTERS_reg_23_45_inst : DFF_X1 port map( D => n3013, CK => n800, Q => 
                           REGISTERS_23_45_port, QN => n_2494);
   REGISTERS_reg_23_44_inst : DFF_X1 port map( D => n3012, CK => n800, Q => 
                           REGISTERS_23_44_port, QN => n_2495);
   REGISTERS_reg_23_43_inst : DFF_X1 port map( D => n3011, CK => n800, Q => 
                           REGISTERS_23_43_port, QN => n_2496);
   REGISTERS_reg_23_42_inst : DFF_X1 port map( D => n3010, CK => n800, Q => 
                           REGISTERS_23_42_port, QN => n_2497);
   REGISTERS_reg_23_41_inst : DFF_X1 port map( D => n3009, CK => n800, Q => 
                           REGISTERS_23_41_port, QN => n_2498);
   REGISTERS_reg_23_40_inst : DFF_X1 port map( D => n3008, CK => n801, Q => 
                           REGISTERS_23_40_port, QN => n_2499);
   REGISTERS_reg_23_39_inst : DFF_X1 port map( D => n3007, CK => n801, Q => 
                           REGISTERS_23_39_port, QN => n_2500);
   REGISTERS_reg_23_38_inst : DFF_X1 port map( D => n3006, CK => n801, Q => 
                           REGISTERS_23_38_port, QN => n_2501);
   REGISTERS_reg_23_37_inst : DFF_X1 port map( D => n3005, CK => n801, Q => 
                           REGISTERS_23_37_port, QN => n_2502);
   REGISTERS_reg_23_36_inst : DFF_X1 port map( D => n3004, CK => n801, Q => 
                           REGISTERS_23_36_port, QN => n_2503);
   REGISTERS_reg_23_35_inst : DFF_X1 port map( D => n3003, CK => n801, Q => 
                           REGISTERS_23_35_port, QN => n_2504);
   REGISTERS_reg_23_34_inst : DFF_X1 port map( D => n3002, CK => n801, Q => 
                           REGISTERS_23_34_port, QN => n_2505);
   REGISTERS_reg_23_33_inst : DFF_X1 port map( D => n3001, CK => n801, Q => 
                           REGISTERS_23_33_port, QN => n_2506);
   REGISTERS_reg_23_32_inst : DFF_X1 port map( D => n3000, CK => n801, Q => 
                           REGISTERS_23_32_port, QN => n_2507);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n2999, CK => n801, Q => 
                           REGISTERS_23_31_port, QN => n_2508);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n2998, CK => n801, Q => 
                           REGISTERS_23_30_port, QN => n_2509);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n2997, CK => n802, Q => 
                           REGISTERS_23_29_port, QN => n_2510);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n2996, CK => n802, Q => 
                           REGISTERS_23_28_port, QN => n_2511);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n2995, CK => n802, Q => 
                           REGISTERS_23_27_port, QN => n_2512);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n2994, CK => n802, Q => 
                           REGISTERS_23_26_port, QN => n_2513);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n2993, CK => n802, Q => 
                           REGISTERS_23_25_port, QN => n_2514);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n2992, CK => n802, Q => 
                           REGISTERS_23_24_port, QN => n_2515);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n2991, CK => n802, Q => 
                           REGISTERS_23_23_port, QN => n_2516);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n2990, CK => n802, Q => 
                           REGISTERS_23_22_port, QN => n_2517);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n2989, CK => n802, Q => 
                           REGISTERS_23_21_port, QN => n_2518);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n2988, CK => n802, Q => 
                           REGISTERS_23_20_port, QN => n_2519);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n2987, CK => n802, Q => 
                           REGISTERS_23_19_port, QN => n_2520);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n2986, CK => n803, Q => 
                           REGISTERS_23_18_port, QN => n_2521);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n2985, CK => n803, Q => 
                           REGISTERS_23_17_port, QN => n_2522);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n2984, CK => n803, Q => 
                           REGISTERS_23_16_port, QN => n_2523);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n2983, CK => n803, Q => 
                           REGISTERS_23_15_port, QN => n_2524);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n2982, CK => n803, Q => 
                           REGISTERS_23_14_port, QN => n_2525);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n2981, CK => n803, Q => 
                           REGISTERS_23_13_port, QN => n_2526);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n2980, CK => n803, Q => 
                           REGISTERS_23_12_port, QN => n_2527);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n2979, CK => n803, Q => 
                           REGISTERS_23_11_port, QN => n_2528);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n2978, CK => n803, Q => 
                           REGISTERS_23_10_port, QN => n_2529);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n2977, CK => n803, Q => 
                           REGISTERS_23_9_port, QN => n_2530);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n2976, CK => n803, Q => 
                           REGISTERS_23_8_port, QN => n_2531);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n2975, CK => n804, Q => 
                           REGISTERS_23_7_port, QN => n_2532);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n2974, CK => n804, Q => 
                           REGISTERS_23_6_port, QN => n_2533);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n2973, CK => n804, Q => 
                           REGISTERS_23_5_port, QN => n_2534);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n2972, CK => n804, Q => 
                           REGISTERS_23_4_port, QN => n_2535);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n2971, CK => n804, Q => 
                           REGISTERS_23_3_port, QN => n_2536);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n2970, CK => n804, Q => 
                           REGISTERS_23_2_port, QN => n_2537);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n2969, CK => n804, Q => 
                           REGISTERS_23_1_port, QN => n_2538);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n2968, CK => n804, Q => 
                           REGISTERS_23_0_port, QN => n_2539);
   REGISTERS_reg_24_63_inst : DFF_X1 port map( D => n2967, CK => n700, Q => 
                           REGISTERS_24_63_port, QN => n_2540);
   REGISTERS_reg_24_62_inst : DFF_X1 port map( D => n2966, CK => n700, Q => 
                           REGISTERS_24_62_port, QN => n_2541);
   REGISTERS_reg_24_61_inst : DFF_X1 port map( D => n2965, CK => n700, Q => 
                           REGISTERS_24_61_port, QN => n_2542);
   REGISTERS_reg_24_60_inst : DFF_X1 port map( D => n2964, CK => n701, Q => 
                           REGISTERS_24_60_port, QN => n_2543);
   REGISTERS_reg_24_59_inst : DFF_X1 port map( D => n2963, CK => n701, Q => 
                           REGISTERS_24_59_port, QN => n_2544);
   REGISTERS_reg_24_58_inst : DFF_X1 port map( D => n2962, CK => n701, Q => 
                           REGISTERS_24_58_port, QN => n_2545);
   REGISTERS_reg_24_57_inst : DFF_X1 port map( D => n2961, CK => n701, Q => 
                           REGISTERS_24_57_port, QN => n_2546);
   REGISTERS_reg_24_56_inst : DFF_X1 port map( D => n2960, CK => n702, Q => 
                           REGISTERS_24_56_port, QN => n_2547);
   REGISTERS_reg_24_55_inst : DFF_X1 port map( D => n2959, CK => n702, Q => 
                           REGISTERS_24_55_port, QN => n_2548);
   REGISTERS_reg_24_54_inst : DFF_X1 port map( D => n2958, CK => n702, Q => 
                           REGISTERS_24_54_port, QN => n_2549);
   REGISTERS_reg_24_53_inst : DFF_X1 port map( D => n2957, CK => n702, Q => 
                           REGISTERS_24_53_port, QN => n_2550);
   REGISTERS_reg_24_52_inst : DFF_X1 port map( D => n2956, CK => n703, Q => 
                           REGISTERS_24_52_port, QN => n_2551);
   REGISTERS_reg_24_51_inst : DFF_X1 port map( D => n2955, CK => n703, Q => 
                           REGISTERS_24_51_port, QN => n_2552);
   REGISTERS_reg_24_50_inst : DFF_X1 port map( D => n2954, CK => n703, Q => 
                           REGISTERS_24_50_port, QN => n_2553);
   REGISTERS_reg_24_49_inst : DFF_X1 port map( D => n2953, CK => n704, Q => 
                           REGISTERS_24_49_port, QN => n_2554);
   REGISTERS_reg_24_48_inst : DFF_X1 port map( D => n2952, CK => n704, Q => 
                           REGISTERS_24_48_port, QN => n_2555);
   REGISTERS_reg_24_47_inst : DFF_X1 port map( D => n2951, CK => n704, Q => 
                           REGISTERS_24_47_port, QN => n_2556);
   REGISTERS_reg_24_46_inst : DFF_X1 port map( D => n2950, CK => n704, Q => 
                           REGISTERS_24_46_port, QN => n_2557);
   REGISTERS_reg_24_45_inst : DFF_X1 port map( D => n2949, CK => n705, Q => 
                           REGISTERS_24_45_port, QN => n_2558);
   REGISTERS_reg_24_44_inst : DFF_X1 port map( D => n2948, CK => n705, Q => 
                           REGISTERS_24_44_port, QN => n_2559);
   REGISTERS_reg_24_43_inst : DFF_X1 port map( D => n2947, CK => n705, Q => 
                           REGISTERS_24_43_port, QN => n_2560);
   REGISTERS_reg_24_42_inst : DFF_X1 port map( D => n2946, CK => n705, Q => 
                           REGISTERS_24_42_port, QN => n_2561);
   REGISTERS_reg_24_41_inst : DFF_X1 port map( D => n2945, CK => n706, Q => 
                           REGISTERS_24_41_port, QN => n_2562);
   REGISTERS_reg_24_40_inst : DFF_X1 port map( D => n2944, CK => n706, Q => 
                           REGISTERS_24_40_port, QN => n_2563);
   REGISTERS_reg_24_39_inst : DFF_X1 port map( D => n2943, CK => n706, Q => 
                           REGISTERS_24_39_port, QN => n_2564);
   REGISTERS_reg_24_38_inst : DFF_X1 port map( D => n2942, CK => n707, Q => 
                           REGISTERS_24_38_port, QN => n_2565);
   REGISTERS_reg_24_37_inst : DFF_X1 port map( D => n2941, CK => n707, Q => 
                           REGISTERS_24_37_port, QN => n_2566);
   REGISTERS_reg_24_36_inst : DFF_X1 port map( D => n2940, CK => n707, Q => 
                           REGISTERS_24_36_port, QN => n_2567);
   REGISTERS_reg_24_35_inst : DFF_X1 port map( D => n2939, CK => n707, Q => 
                           REGISTERS_24_35_port, QN => n_2568);
   REGISTERS_reg_24_34_inst : DFF_X1 port map( D => n2938, CK => n708, Q => 
                           REGISTERS_24_34_port, QN => n_2569);
   REGISTERS_reg_24_33_inst : DFF_X1 port map( D => n2937, CK => n708, Q => 
                           REGISTERS_24_33_port, QN => n_2570);
   REGISTERS_reg_24_32_inst : DFF_X1 port map( D => n2936, CK => n708, Q => 
                           REGISTERS_24_32_port, QN => n_2571);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n2935, CK => n708, Q => 
                           REGISTERS_24_31_port, QN => n_2572);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n2934, CK => n709, Q => 
                           REGISTERS_24_30_port, QN => n_2573);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n2933, CK => n709, Q => 
                           REGISTERS_24_29_port, QN => n_2574);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n2932, CK => n709, Q => 
                           REGISTERS_24_28_port, QN => n_2575);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n2931, CK => n710, Q => 
                           REGISTERS_24_27_port, QN => n_2576);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n2930, CK => n710, Q => 
                           REGISTERS_24_26_port, QN => n_2577);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n2929, CK => n710, Q => 
                           REGISTERS_24_25_port, QN => n_2578);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n2928, CK => n710, Q => 
                           REGISTERS_24_24_port, QN => n_2579);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n2927, CK => n711, Q => 
                           REGISTERS_24_23_port, QN => n_2580);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n2926, CK => n711, Q => 
                           REGISTERS_24_22_port, QN => n_2581);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n2925, CK => n711, Q => 
                           REGISTERS_24_21_port, QN => n_2582);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n2924, CK => n711, Q => 
                           REGISTERS_24_20_port, QN => n_2583);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n2923, CK => n712, Q => 
                           REGISTERS_24_19_port, QN => n_2584);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n2922, CK => n712, Q => 
                           REGISTERS_24_18_port, QN => n_2585);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n2921, CK => n712, Q => 
                           REGISTERS_24_17_port, QN => n_2586);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n2920, CK => n713, Q => 
                           REGISTERS_24_16_port, QN => n_2587);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n2919, CK => n713, Q => 
                           REGISTERS_24_15_port, QN => n_2588);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n2918, CK => n713, Q => 
                           REGISTERS_24_14_port, QN => n_2589);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n2917, CK => n713, Q => 
                           REGISTERS_24_13_port, QN => n_2590);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n2916, CK => n714, Q => 
                           REGISTERS_24_12_port, QN => n_2591);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n2915, CK => n714, Q => 
                           REGISTERS_24_11_port, QN => n_2592);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n2914, CK => n714, Q => 
                           REGISTERS_24_10_port, QN => n_2593);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n2913, CK => n714, Q => 
                           REGISTERS_24_9_port, QN => n_2594);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n2912, CK => n715, Q => 
                           REGISTERS_24_8_port, QN => n_2595);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n2911, CK => n715, Q => 
                           REGISTERS_24_7_port, QN => n_2596);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n2910, CK => n715, Q => 
                           REGISTERS_24_6_port, QN => n_2597);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n2909, CK => n716, Q => 
                           REGISTERS_24_5_port, QN => n_2598);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n2908, CK => n716, Q => 
                           REGISTERS_24_4_port, QN => n_2599);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n2907, CK => n716, Q => 
                           REGISTERS_24_3_port, QN => n_2600);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n2906, CK => n716, Q => 
                           REGISTERS_24_2_port, QN => n_2601);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n2905, CK => n717, Q => 
                           REGISTERS_24_1_port, QN => n_2602);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n2904, CK => n717, Q => 
                           REGISTERS_24_0_port, QN => n_2603);
   REGISTERS_reg_25_63_inst : DFF_X1 port map( D => n2903, CK => n717, Q => 
                           REGISTERS_25_63_port, QN => n_2604);
   REGISTERS_reg_25_62_inst : DFF_X1 port map( D => n2902, CK => n717, Q => 
                           REGISTERS_25_62_port, QN => n_2605);
   REGISTERS_reg_25_61_inst : DFF_X1 port map( D => n2901, CK => n717, Q => 
                           REGISTERS_25_61_port, QN => n_2606);
   REGISTERS_reg_25_60_inst : DFF_X1 port map( D => n2900, CK => n717, Q => 
                           REGISTERS_25_60_port, QN => n_2607);
   REGISTERS_reg_25_59_inst : DFF_X1 port map( D => n2899, CK => n717, Q => 
                           REGISTERS_25_59_port, QN => n_2608);
   REGISTERS_reg_25_58_inst : DFF_X1 port map( D => n2898, CK => n717, Q => 
                           REGISTERS_25_58_port, QN => n_2609);
   REGISTERS_reg_25_57_inst : DFF_X1 port map( D => n2897, CK => n718, Q => 
                           REGISTERS_25_57_port, QN => n_2610);
   REGISTERS_reg_25_56_inst : DFF_X1 port map( D => n2896, CK => n718, Q => 
                           REGISTERS_25_56_port, QN => n_2611);
   REGISTERS_reg_25_55_inst : DFF_X1 port map( D => n2895, CK => n718, Q => 
                           REGISTERS_25_55_port, QN => n_2612);
   REGISTERS_reg_25_54_inst : DFF_X1 port map( D => n2894, CK => n718, Q => 
                           REGISTERS_25_54_port, QN => n_2613);
   REGISTERS_reg_25_53_inst : DFF_X1 port map( D => n2893, CK => n718, Q => 
                           REGISTERS_25_53_port, QN => n_2614);
   REGISTERS_reg_25_52_inst : DFF_X1 port map( D => n2892, CK => n718, Q => 
                           REGISTERS_25_52_port, QN => n_2615);
   REGISTERS_reg_25_51_inst : DFF_X1 port map( D => n2891, CK => n718, Q => 
                           REGISTERS_25_51_port, QN => n_2616);
   REGISTERS_reg_25_50_inst : DFF_X1 port map( D => n2890, CK => n718, Q => 
                           REGISTERS_25_50_port, QN => n_2617);
   REGISTERS_reg_25_49_inst : DFF_X1 port map( D => n2889, CK => n718, Q => 
                           REGISTERS_25_49_port, QN => n_2618);
   REGISTERS_reg_25_48_inst : DFF_X1 port map( D => n2888, CK => n718, Q => 
                           REGISTERS_25_48_port, QN => n_2619);
   REGISTERS_reg_25_47_inst : DFF_X1 port map( D => n2887, CK => n718, Q => 
                           REGISTERS_25_47_port, QN => n_2620);
   REGISTERS_reg_25_46_inst : DFF_X1 port map( D => n2886, CK => n719, Q => 
                           REGISTERS_25_46_port, QN => n_2621);
   REGISTERS_reg_25_45_inst : DFF_X1 port map( D => n2885, CK => n719, Q => 
                           REGISTERS_25_45_port, QN => n_2622);
   REGISTERS_reg_25_44_inst : DFF_X1 port map( D => n2884, CK => n719, Q => 
                           REGISTERS_25_44_port, QN => n_2623);
   REGISTERS_reg_25_43_inst : DFF_X1 port map( D => n2883, CK => n719, Q => 
                           REGISTERS_25_43_port, QN => n_2624);
   REGISTERS_reg_25_42_inst : DFF_X1 port map( D => n2882, CK => n719, Q => 
                           REGISTERS_25_42_port, QN => n_2625);
   REGISTERS_reg_25_41_inst : DFF_X1 port map( D => n2881, CK => n719, Q => 
                           REGISTERS_25_41_port, QN => n_2626);
   REGISTERS_reg_25_40_inst : DFF_X1 port map( D => n2880, CK => n719, Q => 
                           REGISTERS_25_40_port, QN => n_2627);
   REGISTERS_reg_25_39_inst : DFF_X1 port map( D => n2879, CK => n719, Q => 
                           REGISTERS_25_39_port, QN => n_2628);
   REGISTERS_reg_25_38_inst : DFF_X1 port map( D => n2878, CK => n719, Q => 
                           REGISTERS_25_38_port, QN => n_2629);
   REGISTERS_reg_25_37_inst : DFF_X1 port map( D => n2877, CK => n719, Q => 
                           REGISTERS_25_37_port, QN => n_2630);
   REGISTERS_reg_25_36_inst : DFF_X1 port map( D => n2876, CK => n719, Q => 
                           REGISTERS_25_36_port, QN => n_2631);
   REGISTERS_reg_25_35_inst : DFF_X1 port map( D => n2875, CK => n720, Q => 
                           REGISTERS_25_35_port, QN => n_2632);
   REGISTERS_reg_25_34_inst : DFF_X1 port map( D => n2874, CK => n720, Q => 
                           REGISTERS_25_34_port, QN => n_2633);
   REGISTERS_reg_25_33_inst : DFF_X1 port map( D => n2873, CK => n720, Q => 
                           REGISTERS_25_33_port, QN => n_2634);
   REGISTERS_reg_25_32_inst : DFF_X1 port map( D => n2872, CK => n720, Q => 
                           REGISTERS_25_32_port, QN => n_2635);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n2871, CK => n720, Q => 
                           REGISTERS_25_31_port, QN => n_2636);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n2870, CK => n720, Q => 
                           REGISTERS_25_30_port, QN => n_2637);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n2869, CK => n720, Q => 
                           REGISTERS_25_29_port, QN => n_2638);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n2868, CK => n720, Q => 
                           REGISTERS_25_28_port, QN => n_2639);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n2867, CK => n720, Q => 
                           REGISTERS_25_27_port, QN => n_2640);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n2866, CK => n720, Q => 
                           REGISTERS_25_26_port, QN => n_2641);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n2865, CK => n720, Q => 
                           REGISTERS_25_25_port, QN => n_2642);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n2864, CK => n721, Q => 
                           REGISTERS_25_24_port, QN => n_2643);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n2863, CK => n721, Q => 
                           REGISTERS_25_23_port, QN => n_2644);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n2862, CK => n721, Q => 
                           REGISTERS_25_22_port, QN => n_2645);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n2861, CK => n721, Q => 
                           REGISTERS_25_21_port, QN => n_2646);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n2860, CK => n721, Q => 
                           REGISTERS_25_20_port, QN => n_2647);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n2859, CK => n721, Q => 
                           REGISTERS_25_19_port, QN => n_2648);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n2858, CK => n721, Q => 
                           REGISTERS_25_18_port, QN => n_2649);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n2857, CK => n721, Q => 
                           REGISTERS_25_17_port, QN => n_2650);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n2856, CK => n721, Q => 
                           REGISTERS_25_16_port, QN => n_2651);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n2855, CK => n721, Q => 
                           REGISTERS_25_15_port, QN => n_2652);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n2854, CK => n721, Q => 
                           REGISTERS_25_14_port, QN => n_2653);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n2853, CK => n722, Q => 
                           REGISTERS_25_13_port, QN => n_2654);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n2852, CK => n722, Q => 
                           REGISTERS_25_12_port, QN => n_2655);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n2851, CK => n722, Q => 
                           REGISTERS_25_11_port, QN => n_2656);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n2850, CK => n722, Q => 
                           REGISTERS_25_10_port, QN => n_2657);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n2849, CK => n722, Q => 
                           REGISTERS_25_9_port, QN => n_2658);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n2848, CK => n722, Q => 
                           REGISTERS_25_8_port, QN => n_2659);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n2847, CK => n722, Q => 
                           REGISTERS_25_7_port, QN => n_2660);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n2846, CK => n722, Q => 
                           REGISTERS_25_6_port, QN => n_2661);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n2845, CK => n722, Q => 
                           REGISTERS_25_5_port, QN => n_2662);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n2844, CK => n722, Q => 
                           REGISTERS_25_4_port, QN => n_2663);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n2843, CK => n722, Q => 
                           REGISTERS_25_3_port, QN => n_2664);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n2842, CK => n723, Q => 
                           REGISTERS_25_2_port, QN => n_2665);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n2841, CK => n723, Q => 
                           REGISTERS_25_1_port, QN => n_2666);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n2840, CK => n723, Q => 
                           REGISTERS_25_0_port, QN => n_2667);
   REGISTERS_reg_26_63_inst : DFF_X1 port map( D => n2839, CK => n723, Q => 
                           REGISTERS_26_63_port, QN => n_2668);
   REGISTERS_reg_26_62_inst : DFF_X1 port map( D => n2838, CK => n723, Q => 
                           REGISTERS_26_62_port, QN => n_2669);
   REGISTERS_reg_26_61_inst : DFF_X1 port map( D => n2837, CK => n723, Q => 
                           REGISTERS_26_61_port, QN => n_2670);
   REGISTERS_reg_26_60_inst : DFF_X1 port map( D => n2836, CK => n723, Q => 
                           REGISTERS_26_60_port, QN => n_2671);
   REGISTERS_reg_26_59_inst : DFF_X1 port map( D => n2835, CK => n723, Q => 
                           REGISTERS_26_59_port, QN => n_2672);
   REGISTERS_reg_26_58_inst : DFF_X1 port map( D => n2834, CK => n723, Q => 
                           REGISTERS_26_58_port, QN => n_2673);
   REGISTERS_reg_26_57_inst : DFF_X1 port map( D => n2833, CK => n723, Q => 
                           REGISTERS_26_57_port, QN => n_2674);
   REGISTERS_reg_26_56_inst : DFF_X1 port map( D => n2832, CK => n723, Q => 
                           REGISTERS_26_56_port, QN => n_2675);
   REGISTERS_reg_26_55_inst : DFF_X1 port map( D => n2831, CK => n724, Q => 
                           REGISTERS_26_55_port, QN => n_2676);
   REGISTERS_reg_26_54_inst : DFF_X1 port map( D => n2830, CK => n724, Q => 
                           REGISTERS_26_54_port, QN => n_2677);
   REGISTERS_reg_26_53_inst : DFF_X1 port map( D => n2829, CK => n724, Q => 
                           REGISTERS_26_53_port, QN => n_2678);
   REGISTERS_reg_26_52_inst : DFF_X1 port map( D => n2828, CK => n724, Q => 
                           REGISTERS_26_52_port, QN => n_2679);
   REGISTERS_reg_26_51_inst : DFF_X1 port map( D => n2827, CK => n724, Q => 
                           REGISTERS_26_51_port, QN => n_2680);
   REGISTERS_reg_26_50_inst : DFF_X1 port map( D => n2826, CK => n724, Q => 
                           REGISTERS_26_50_port, QN => n_2681);
   REGISTERS_reg_26_49_inst : DFF_X1 port map( D => n2825, CK => n724, Q => 
                           REGISTERS_26_49_port, QN => n_2682);
   REGISTERS_reg_26_48_inst : DFF_X1 port map( D => n2824, CK => n724, Q => 
                           REGISTERS_26_48_port, QN => n_2683);
   REGISTERS_reg_26_47_inst : DFF_X1 port map( D => n2823, CK => n724, Q => 
                           REGISTERS_26_47_port, QN => n_2684);
   REGISTERS_reg_26_46_inst : DFF_X1 port map( D => n2822, CK => n724, Q => 
                           REGISTERS_26_46_port, QN => n_2685);
   REGISTERS_reg_26_45_inst : DFF_X1 port map( D => n2821, CK => n724, Q => 
                           REGISTERS_26_45_port, QN => n_2686);
   REGISTERS_reg_26_44_inst : DFF_X1 port map( D => n2820, CK => n725, Q => 
                           REGISTERS_26_44_port, QN => n_2687);
   REGISTERS_reg_26_43_inst : DFF_X1 port map( D => n2819, CK => n725, Q => 
                           REGISTERS_26_43_port, QN => n_2688);
   REGISTERS_reg_26_42_inst : DFF_X1 port map( D => n2818, CK => n725, Q => 
                           REGISTERS_26_42_port, QN => n_2689);
   REGISTERS_reg_26_41_inst : DFF_X1 port map( D => n2817, CK => n725, Q => 
                           REGISTERS_26_41_port, QN => n_2690);
   REGISTERS_reg_26_40_inst : DFF_X1 port map( D => n2816, CK => n725, Q => 
                           REGISTERS_26_40_port, QN => n_2691);
   REGISTERS_reg_26_39_inst : DFF_X1 port map( D => n2815, CK => n725, Q => 
                           REGISTERS_26_39_port, QN => n_2692);
   REGISTERS_reg_26_38_inst : DFF_X1 port map( D => n2814, CK => n725, Q => 
                           REGISTERS_26_38_port, QN => n_2693);
   REGISTERS_reg_26_37_inst : DFF_X1 port map( D => n2813, CK => n725, Q => 
                           REGISTERS_26_37_port, QN => n_2694);
   REGISTERS_reg_26_36_inst : DFF_X1 port map( D => n2812, CK => n725, Q => 
                           REGISTERS_26_36_port, QN => n_2695);
   REGISTERS_reg_26_35_inst : DFF_X1 port map( D => n2811, CK => n725, Q => 
                           REGISTERS_26_35_port, QN => n_2696);
   REGISTERS_reg_26_34_inst : DFF_X1 port map( D => n2810, CK => n725, Q => 
                           REGISTERS_26_34_port, QN => n_2697);
   REGISTERS_reg_26_33_inst : DFF_X1 port map( D => n2809, CK => n726, Q => 
                           REGISTERS_26_33_port, QN => n_2698);
   REGISTERS_reg_26_32_inst : DFF_X1 port map( D => n2808, CK => n726, Q => 
                           REGISTERS_26_32_port, QN => n_2699);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n2807, CK => n726, Q => 
                           REGISTERS_26_31_port, QN => n_2700);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n2806, CK => n726, Q => 
                           REGISTERS_26_30_port, QN => n_2701);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n2805, CK => n726, Q => 
                           REGISTERS_26_29_port, QN => n_2702);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n2804, CK => n726, Q => 
                           REGISTERS_26_28_port, QN => n_2703);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n2803, CK => n726, Q => 
                           REGISTERS_26_27_port, QN => n_2704);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n2802, CK => n726, Q => 
                           REGISTERS_26_26_port, QN => n_2705);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n2801, CK => n726, Q => 
                           REGISTERS_26_25_port, QN => n_2706);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n2800, CK => n726, Q => 
                           REGISTERS_26_24_port, QN => n_2707);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n2799, CK => n726, Q => 
                           REGISTERS_26_23_port, QN => n_2708);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n2798, CK => n727, Q => 
                           REGISTERS_26_22_port, QN => n_2709);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n2797, CK => n727, Q => 
                           REGISTERS_26_21_port, QN => n_2710);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n2796, CK => n727, Q => 
                           REGISTERS_26_20_port, QN => n_2711);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n2795, CK => n727, Q => 
                           REGISTERS_26_19_port, QN => n_2712);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n2794, CK => n727, Q => 
                           REGISTERS_26_18_port, QN => n_2713);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n2793, CK => n727, Q => 
                           REGISTERS_26_17_port, QN => n_2714);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n2792, CK => n727, Q => 
                           REGISTERS_26_16_port, QN => n_2715);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n2791, CK => n727, Q => 
                           REGISTERS_26_15_port, QN => n_2716);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n2790, CK => n727, Q => 
                           REGISTERS_26_14_port, QN => n_2717);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n2789, CK => n727, Q => 
                           REGISTERS_26_13_port, QN => n_2718);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n2788, CK => n727, Q => 
                           REGISTERS_26_12_port, QN => n_2719);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n2787, CK => n728, Q => 
                           REGISTERS_26_11_port, QN => n_2720);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n2786, CK => n728, Q => 
                           REGISTERS_26_10_port, QN => n_2721);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n2785, CK => n728, Q => 
                           REGISTERS_26_9_port, QN => n_2722);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n2784, CK => n728, Q => 
                           REGISTERS_26_8_port, QN => n_2723);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n2783, CK => n728, Q => 
                           REGISTERS_26_7_port, QN => n_2724);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n2782, CK => n728, Q => 
                           REGISTERS_26_6_port, QN => n_2725);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n2781, CK => n728, Q => 
                           REGISTERS_26_5_port, QN => n_2726);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n2780, CK => n728, Q => 
                           REGISTERS_26_4_port, QN => n_2727);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n2779, CK => n728, Q => 
                           REGISTERS_26_3_port, QN => n_2728);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n2778, CK => n728, Q => 
                           REGISTERS_26_2_port, QN => n_2729);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n2777, CK => n728, Q => 
                           REGISTERS_26_1_port, QN => n_2730);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n2776, CK => n729, Q => 
                           REGISTERS_26_0_port, QN => n_2731);
   REGISTERS_reg_27_63_inst : DFF_X1 port map( D => n2775, CK => n729, Q => 
                           REGISTERS_27_63_port, QN => n_2732);
   REGISTERS_reg_27_62_inst : DFF_X1 port map( D => n2774, CK => n729, Q => 
                           REGISTERS_27_62_port, QN => n_2733);
   REGISTERS_reg_27_61_inst : DFF_X1 port map( D => n2773, CK => n729, Q => 
                           REGISTERS_27_61_port, QN => n_2734);
   REGISTERS_reg_27_60_inst : DFF_X1 port map( D => n2772, CK => n729, Q => 
                           REGISTERS_27_60_port, QN => n_2735);
   REGISTERS_reg_27_59_inst : DFF_X1 port map( D => n2771, CK => n729, Q => 
                           REGISTERS_27_59_port, QN => n_2736);
   REGISTERS_reg_27_58_inst : DFF_X1 port map( D => n2770, CK => n729, Q => 
                           REGISTERS_27_58_port, QN => n_2737);
   REGISTERS_reg_27_57_inst : DFF_X1 port map( D => n2769, CK => n729, Q => 
                           REGISTERS_27_57_port, QN => n_2738);
   REGISTERS_reg_27_56_inst : DFF_X1 port map( D => n2768, CK => n729, Q => 
                           REGISTERS_27_56_port, QN => n_2739);
   REGISTERS_reg_27_55_inst : DFF_X1 port map( D => n2767, CK => n729, Q => 
                           REGISTERS_27_55_port, QN => n_2740);
   REGISTERS_reg_27_54_inst : DFF_X1 port map( D => n2766, CK => n729, Q => 
                           REGISTERS_27_54_port, QN => n_2741);
   REGISTERS_reg_27_53_inst : DFF_X1 port map( D => n2765, CK => n730, Q => 
                           REGISTERS_27_53_port, QN => n_2742);
   REGISTERS_reg_27_52_inst : DFF_X1 port map( D => n2764, CK => n730, Q => 
                           REGISTERS_27_52_port, QN => n_2743);
   REGISTERS_reg_27_51_inst : DFF_X1 port map( D => n2763, CK => n730, Q => 
                           REGISTERS_27_51_port, QN => n_2744);
   REGISTERS_reg_27_50_inst : DFF_X1 port map( D => n2762, CK => n730, Q => 
                           REGISTERS_27_50_port, QN => n_2745);
   REGISTERS_reg_27_49_inst : DFF_X1 port map( D => n2761, CK => n730, Q => 
                           REGISTERS_27_49_port, QN => n_2746);
   REGISTERS_reg_27_48_inst : DFF_X1 port map( D => n2760, CK => n730, Q => 
                           REGISTERS_27_48_port, QN => n_2747);
   REGISTERS_reg_27_47_inst : DFF_X1 port map( D => n2759, CK => n730, Q => 
                           REGISTERS_27_47_port, QN => n_2748);
   REGISTERS_reg_27_46_inst : DFF_X1 port map( D => n2758, CK => n730, Q => 
                           REGISTERS_27_46_port, QN => n_2749);
   REGISTERS_reg_27_45_inst : DFF_X1 port map( D => n2757, CK => n730, Q => 
                           REGISTERS_27_45_port, QN => n_2750);
   REGISTERS_reg_27_44_inst : DFF_X1 port map( D => n2756, CK => n730, Q => 
                           REGISTERS_27_44_port, QN => n_2751);
   REGISTERS_reg_27_43_inst : DFF_X1 port map( D => n2755, CK => n730, Q => 
                           REGISTERS_27_43_port, QN => n_2752);
   REGISTERS_reg_27_42_inst : DFF_X1 port map( D => n2754, CK => n731, Q => 
                           REGISTERS_27_42_port, QN => n_2753);
   REGISTERS_reg_27_41_inst : DFF_X1 port map( D => n2753, CK => n731, Q => 
                           REGISTERS_27_41_port, QN => n_2754);
   REGISTERS_reg_27_40_inst : DFF_X1 port map( D => n2752, CK => n731, Q => 
                           REGISTERS_27_40_port, QN => n_2755);
   REGISTERS_reg_27_39_inst : DFF_X1 port map( D => n2751, CK => n731, Q => 
                           REGISTERS_27_39_port, QN => n_2756);
   REGISTERS_reg_27_38_inst : DFF_X1 port map( D => n2750, CK => n731, Q => 
                           REGISTERS_27_38_port, QN => n_2757);
   REGISTERS_reg_27_37_inst : DFF_X1 port map( D => n2749, CK => n731, Q => 
                           REGISTERS_27_37_port, QN => n_2758);
   REGISTERS_reg_27_36_inst : DFF_X1 port map( D => n2748, CK => n731, Q => 
                           REGISTERS_27_36_port, QN => n_2759);
   REGISTERS_reg_27_35_inst : DFF_X1 port map( D => n2747, CK => n731, Q => 
                           REGISTERS_27_35_port, QN => n_2760);
   REGISTERS_reg_27_34_inst : DFF_X1 port map( D => n2746, CK => n731, Q => 
                           REGISTERS_27_34_port, QN => n_2761);
   REGISTERS_reg_27_33_inst : DFF_X1 port map( D => n2745, CK => n731, Q => 
                           REGISTERS_27_33_port, QN => n_2762);
   REGISTERS_reg_27_32_inst : DFF_X1 port map( D => n2744, CK => n731, Q => 
                           REGISTERS_27_32_port, QN => n_2763);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n2743, CK => n732, Q => 
                           REGISTERS_27_31_port, QN => n_2764);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n2742, CK => n732, Q => 
                           REGISTERS_27_30_port, QN => n_2765);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n2741, CK => n732, Q => 
                           REGISTERS_27_29_port, QN => n_2766);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n2740, CK => n732, Q => 
                           REGISTERS_27_28_port, QN => n_2767);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n2739, CK => n732, Q => 
                           REGISTERS_27_27_port, QN => n_2768);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n2738, CK => n732, Q => 
                           REGISTERS_27_26_port, QN => n_2769);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n2737, CK => n732, Q => 
                           REGISTERS_27_25_port, QN => n_2770);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n2736, CK => n732, Q => 
                           REGISTERS_27_24_port, QN => n_2771);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n2735, CK => n732, Q => 
                           REGISTERS_27_23_port, QN => n_2772);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n2734, CK => n732, Q => 
                           REGISTERS_27_22_port, QN => n_2773);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n2733, CK => n732, Q => 
                           REGISTERS_27_21_port, QN => n_2774);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n2732, CK => n733, Q => 
                           REGISTERS_27_20_port, QN => n_2775);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n2731, CK => n733, Q => 
                           REGISTERS_27_19_port, QN => n_2776);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n2730, CK => n733, Q => 
                           REGISTERS_27_18_port, QN => n_2777);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n2729, CK => n733, Q => 
                           REGISTERS_27_17_port, QN => n_2778);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n2728, CK => n733, Q => 
                           REGISTERS_27_16_port, QN => n_2779);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n2727, CK => n733, Q => 
                           REGISTERS_27_15_port, QN => n_2780);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n2726, CK => n733, Q => 
                           REGISTERS_27_14_port, QN => n_2781);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n2725, CK => n733, Q => 
                           REGISTERS_27_13_port, QN => n_2782);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n2724, CK => n733, Q => 
                           REGISTERS_27_12_port, QN => n_2783);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n2723, CK => n733, Q => 
                           REGISTERS_27_11_port, QN => n_2784);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n2722, CK => n733, Q => 
                           REGISTERS_27_10_port, QN => n_2785);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n2721, CK => n734, Q => 
                           REGISTERS_27_9_port, QN => n_2786);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n2720, CK => n734, Q => 
                           REGISTERS_27_8_port, QN => n_2787);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n2719, CK => n734, Q => 
                           REGISTERS_27_7_port, QN => n_2788);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n2718, CK => n734, Q => 
                           REGISTERS_27_6_port, QN => n_2789);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n2717, CK => n734, Q => 
                           REGISTERS_27_5_port, QN => n_2790);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n2716, CK => n734, Q => 
                           REGISTERS_27_4_port, QN => n_2791);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n2715, CK => n734, Q => 
                           REGISTERS_27_3_port, QN => n_2792);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n2714, CK => n734, Q => 
                           REGISTERS_27_2_port, QN => n_2793);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n2713, CK => n734, Q => 
                           REGISTERS_27_1_port, QN => n_2794);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n2712, CK => n734, Q => 
                           REGISTERS_27_0_port, QN => n_2795);
   REGISTERS_reg_28_63_inst : DFF_X1 port map( D => n2711, CK => n734, Q => 
                           REGISTERS_28_63_port, QN => n_2796);
   REGISTERS_reg_28_62_inst : DFF_X1 port map( D => n2710, CK => n735, Q => 
                           REGISTERS_28_62_port, QN => n_2797);
   REGISTERS_reg_28_61_inst : DFF_X1 port map( D => n2709, CK => n735, Q => 
                           REGISTERS_28_61_port, QN => n_2798);
   REGISTERS_reg_28_60_inst : DFF_X1 port map( D => n2708, CK => n735, Q => 
                           REGISTERS_28_60_port, QN => n_2799);
   REGISTERS_reg_28_59_inst : DFF_X1 port map( D => n2707, CK => n735, Q => 
                           REGISTERS_28_59_port, QN => n_2800);
   REGISTERS_reg_28_58_inst : DFF_X1 port map( D => n2706, CK => n735, Q => 
                           REGISTERS_28_58_port, QN => n_2801);
   REGISTERS_reg_28_57_inst : DFF_X1 port map( D => n2705, CK => n735, Q => 
                           REGISTERS_28_57_port, QN => n_2802);
   REGISTERS_reg_28_56_inst : DFF_X1 port map( D => n2704, CK => n735, Q => 
                           REGISTERS_28_56_port, QN => n_2803);
   REGISTERS_reg_28_55_inst : DFF_X1 port map( D => n2703, CK => n735, Q => 
                           REGISTERS_28_55_port, QN => n_2804);
   REGISTERS_reg_28_54_inst : DFF_X1 port map( D => n2702, CK => n735, Q => 
                           REGISTERS_28_54_port, QN => n_2805);
   REGISTERS_reg_28_53_inst : DFF_X1 port map( D => n2701, CK => n735, Q => 
                           REGISTERS_28_53_port, QN => n_2806);
   REGISTERS_reg_28_52_inst : DFF_X1 port map( D => n2700, CK => n735, Q => 
                           REGISTERS_28_52_port, QN => n_2807);
   REGISTERS_reg_28_51_inst : DFF_X1 port map( D => n2699, CK => n736, Q => 
                           REGISTERS_28_51_port, QN => n_2808);
   REGISTERS_reg_28_50_inst : DFF_X1 port map( D => n2698, CK => n736, Q => 
                           REGISTERS_28_50_port, QN => n_2809);
   REGISTERS_reg_28_49_inst : DFF_X1 port map( D => n2697, CK => n736, Q => 
                           REGISTERS_28_49_port, QN => n_2810);
   REGISTERS_reg_28_48_inst : DFF_X1 port map( D => n2696, CK => n736, Q => 
                           REGISTERS_28_48_port, QN => n_2811);
   REGISTERS_reg_28_47_inst : DFF_X1 port map( D => n2695, CK => n736, Q => 
                           REGISTERS_28_47_port, QN => n_2812);
   REGISTERS_reg_28_46_inst : DFF_X1 port map( D => n2694, CK => n736, Q => 
                           REGISTERS_28_46_port, QN => n_2813);
   REGISTERS_reg_28_45_inst : DFF_X1 port map( D => n2693, CK => n736, Q => 
                           REGISTERS_28_45_port, QN => n_2814);
   REGISTERS_reg_28_44_inst : DFF_X1 port map( D => n2692, CK => n736, Q => 
                           REGISTERS_28_44_port, QN => n_2815);
   REGISTERS_reg_28_43_inst : DFF_X1 port map( D => n2691, CK => n736, Q => 
                           REGISTERS_28_43_port, QN => n_2816);
   REGISTERS_reg_28_42_inst : DFF_X1 port map( D => n2690, CK => n736, Q => 
                           REGISTERS_28_42_port, QN => n_2817);
   REGISTERS_reg_28_41_inst : DFF_X1 port map( D => n2689, CK => n736, Q => 
                           REGISTERS_28_41_port, QN => n_2818);
   REGISTERS_reg_28_40_inst : DFF_X1 port map( D => n2688, CK => n737, Q => 
                           REGISTERS_28_40_port, QN => n_2819);
   REGISTERS_reg_28_39_inst : DFF_X1 port map( D => n2687, CK => n737, Q => 
                           REGISTERS_28_39_port, QN => n_2820);
   REGISTERS_reg_28_38_inst : DFF_X1 port map( D => n2686, CK => n737, Q => 
                           REGISTERS_28_38_port, QN => n_2821);
   REGISTERS_reg_28_37_inst : DFF_X1 port map( D => n2685, CK => n737, Q => 
                           REGISTERS_28_37_port, QN => n_2822);
   REGISTERS_reg_28_36_inst : DFF_X1 port map( D => n2684, CK => n737, Q => 
                           REGISTERS_28_36_port, QN => n_2823);
   REGISTERS_reg_28_35_inst : DFF_X1 port map( D => n2683, CK => n737, Q => 
                           REGISTERS_28_35_port, QN => n_2824);
   REGISTERS_reg_28_34_inst : DFF_X1 port map( D => n2682, CK => n737, Q => 
                           REGISTERS_28_34_port, QN => n_2825);
   REGISTERS_reg_28_33_inst : DFF_X1 port map( D => n2681, CK => n737, Q => 
                           REGISTERS_28_33_port, QN => n_2826);
   REGISTERS_reg_28_32_inst : DFF_X1 port map( D => n2680, CK => n737, Q => 
                           REGISTERS_28_32_port, QN => n_2827);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n2679, CK => n737, Q => 
                           REGISTERS_28_31_port, QN => n_2828);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n2678, CK => n737, Q => 
                           REGISTERS_28_30_port, QN => n_2829);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n2677, CK => n738, Q => 
                           REGISTERS_28_29_port, QN => n_2830);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n2676, CK => n738, Q => 
                           REGISTERS_28_28_port, QN => n_2831);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n2675, CK => n738, Q => 
                           REGISTERS_28_27_port, QN => n_2832);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n2674, CK => n738, Q => 
                           REGISTERS_28_26_port, QN => n_2833);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n2673, CK => n738, Q => 
                           REGISTERS_28_25_port, QN => n_2834);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n2672, CK => n738, Q => 
                           REGISTERS_28_24_port, QN => n_2835);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n2671, CK => n738, Q => 
                           REGISTERS_28_23_port, QN => n_2836);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n2670, CK => n738, Q => 
                           REGISTERS_28_22_port, QN => n_2837);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n2669, CK => n738, Q => 
                           REGISTERS_28_21_port, QN => n_2838);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n2668, CK => n738, Q => 
                           REGISTERS_28_20_port, QN => n_2839);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n2667, CK => n738, Q => 
                           REGISTERS_28_19_port, QN => n_2840);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n2666, CK => n739, Q => 
                           REGISTERS_28_18_port, QN => n_2841);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n2665, CK => n739, Q => 
                           REGISTERS_28_17_port, QN => n_2842);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n2664, CK => n739, Q => 
                           REGISTERS_28_16_port, QN => n_2843);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n2663, CK => n739, Q => 
                           REGISTERS_28_15_port, QN => n_2844);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n2662, CK => n739, Q => 
                           REGISTERS_28_14_port, QN => n_2845);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n2661, CK => n739, Q => 
                           REGISTERS_28_13_port, QN => n_2846);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n2660, CK => n739, Q => 
                           REGISTERS_28_12_port, QN => n_2847);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n2659, CK => n739, Q => 
                           REGISTERS_28_11_port, QN => n_2848);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n2658, CK => n739, Q => 
                           REGISTERS_28_10_port, QN => n_2849);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n2657, CK => n739, Q => 
                           REGISTERS_28_9_port, QN => n_2850);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n2656, CK => n739, Q => 
                           REGISTERS_28_8_port, QN => n_2851);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n2655, CK => n740, Q => 
                           REGISTERS_28_7_port, QN => n_2852);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n2654, CK => n740, Q => 
                           REGISTERS_28_6_port, QN => n_2853);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n2653, CK => n740, Q => 
                           REGISTERS_28_5_port, QN => n_2854);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n2652, CK => n740, Q => 
                           REGISTERS_28_4_port, QN => n_2855);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n2651, CK => n740, Q => 
                           REGISTERS_28_3_port, QN => n_2856);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n2650, CK => n740, Q => 
                           REGISTERS_28_2_port, QN => n_2857);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n2649, CK => n740, Q => 
                           REGISTERS_28_1_port, QN => n_2858);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n2648, CK => n740, Q => 
                           REGISTERS_28_0_port, QN => n_2859);
   REGISTERS_reg_29_63_inst : DFF_X1 port map( D => n2647, CK => n740, Q => 
                           REGISTERS_29_63_port, QN => n_2860);
   REGISTERS_reg_29_62_inst : DFF_X1 port map( D => n2646, CK => n740, Q => 
                           REGISTERS_29_62_port, QN => n_2861);
   REGISTERS_reg_29_61_inst : DFF_X1 port map( D => n2645, CK => n740, Q => 
                           REGISTERS_29_61_port, QN => n_2862);
   REGISTERS_reg_29_60_inst : DFF_X1 port map( D => n2644, CK => n741, Q => 
                           REGISTERS_29_60_port, QN => n_2863);
   REGISTERS_reg_29_59_inst : DFF_X1 port map( D => n2643, CK => n741, Q => 
                           REGISTERS_29_59_port, QN => n_2864);
   REGISTERS_reg_29_58_inst : DFF_X1 port map( D => n2642, CK => n741, Q => 
                           REGISTERS_29_58_port, QN => n_2865);
   REGISTERS_reg_29_57_inst : DFF_X1 port map( D => n2641, CK => n741, Q => 
                           REGISTERS_29_57_port, QN => n_2866);
   REGISTERS_reg_29_56_inst : DFF_X1 port map( D => n2640, CK => n741, Q => 
                           REGISTERS_29_56_port, QN => n_2867);
   REGISTERS_reg_29_55_inst : DFF_X1 port map( D => n2639, CK => n741, Q => 
                           REGISTERS_29_55_port, QN => n_2868);
   REGISTERS_reg_29_54_inst : DFF_X1 port map( D => n2638, CK => n741, Q => 
                           REGISTERS_29_54_port, QN => n_2869);
   REGISTERS_reg_29_53_inst : DFF_X1 port map( D => n2637, CK => n741, Q => 
                           REGISTERS_29_53_port, QN => n_2870);
   REGISTERS_reg_29_52_inst : DFF_X1 port map( D => n2636, CK => n741, Q => 
                           REGISTERS_29_52_port, QN => n_2871);
   REGISTERS_reg_29_51_inst : DFF_X1 port map( D => n2635, CK => n741, Q => 
                           REGISTERS_29_51_port, QN => n_2872);
   REGISTERS_reg_29_50_inst : DFF_X1 port map( D => n2634, CK => n741, Q => 
                           REGISTERS_29_50_port, QN => n_2873);
   REGISTERS_reg_29_49_inst : DFF_X1 port map( D => n2633, CK => n742, Q => 
                           REGISTERS_29_49_port, QN => n_2874);
   REGISTERS_reg_29_48_inst : DFF_X1 port map( D => n2632, CK => n742, Q => 
                           REGISTERS_29_48_port, QN => n_2875);
   REGISTERS_reg_29_47_inst : DFF_X1 port map( D => n2631, CK => n742, Q => 
                           REGISTERS_29_47_port, QN => n_2876);
   REGISTERS_reg_29_46_inst : DFF_X1 port map( D => n2630, CK => n742, Q => 
                           REGISTERS_29_46_port, QN => n_2877);
   REGISTERS_reg_29_45_inst : DFF_X1 port map( D => n2629, CK => n742, Q => 
                           REGISTERS_29_45_port, QN => n_2878);
   REGISTERS_reg_29_44_inst : DFF_X1 port map( D => n2628, CK => n742, Q => 
                           REGISTERS_29_44_port, QN => n_2879);
   REGISTERS_reg_29_43_inst : DFF_X1 port map( D => n2627, CK => n742, Q => 
                           REGISTERS_29_43_port, QN => n_2880);
   REGISTERS_reg_29_42_inst : DFF_X1 port map( D => n2626, CK => n742, Q => 
                           REGISTERS_29_42_port, QN => n_2881);
   REGISTERS_reg_29_41_inst : DFF_X1 port map( D => n2625, CK => n742, Q => 
                           REGISTERS_29_41_port, QN => n_2882);
   REGISTERS_reg_29_40_inst : DFF_X1 port map( D => n2624, CK => n742, Q => 
                           REGISTERS_29_40_port, QN => n_2883);
   REGISTERS_reg_29_39_inst : DFF_X1 port map( D => n2623, CK => n742, Q => 
                           REGISTERS_29_39_port, QN => n_2884);
   REGISTERS_reg_29_38_inst : DFF_X1 port map( D => n2622, CK => n743, Q => 
                           REGISTERS_29_38_port, QN => n_2885);
   REGISTERS_reg_29_37_inst : DFF_X1 port map( D => n2621, CK => n743, Q => 
                           REGISTERS_29_37_port, QN => n_2886);
   REGISTERS_reg_29_36_inst : DFF_X1 port map( D => n2620, CK => n743, Q => 
                           REGISTERS_29_36_port, QN => n_2887);
   REGISTERS_reg_29_35_inst : DFF_X1 port map( D => n2619, CK => n743, Q => 
                           REGISTERS_29_35_port, QN => n_2888);
   REGISTERS_reg_29_34_inst : DFF_X1 port map( D => n2618, CK => n743, Q => 
                           REGISTERS_29_34_port, QN => n_2889);
   REGISTERS_reg_29_33_inst : DFF_X1 port map( D => n2617, CK => n743, Q => 
                           REGISTERS_29_33_port, QN => n_2890);
   REGISTERS_reg_29_32_inst : DFF_X1 port map( D => n2616, CK => n743, Q => 
                           REGISTERS_29_32_port, QN => n_2891);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n2615, CK => n743, Q => 
                           REGISTERS_29_31_port, QN => n_2892);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n2614, CK => n743, Q => 
                           REGISTERS_29_30_port, QN => n_2893);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n2613, CK => n743, Q => 
                           REGISTERS_29_29_port, QN => n_2894);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n2612, CK => n743, Q => 
                           REGISTERS_29_28_port, QN => n_2895);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n2611, CK => n744, Q => 
                           REGISTERS_29_27_port, QN => n_2896);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n2610, CK => n744, Q => 
                           REGISTERS_29_26_port, QN => n_2897);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n2609, CK => n744, Q => 
                           REGISTERS_29_25_port, QN => n_2898);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n2608, CK => n744, Q => 
                           REGISTERS_29_24_port, QN => n_2899);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n2607, CK => n744, Q => 
                           REGISTERS_29_23_port, QN => n_2900);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n2606, CK => n744, Q => 
                           REGISTERS_29_22_port, QN => n_2901);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n2605, CK => n744, Q => 
                           REGISTERS_29_21_port, QN => n_2902);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n2604, CK => n744, Q => 
                           REGISTERS_29_20_port, QN => n_2903);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n2603, CK => n744, Q => 
                           REGISTERS_29_19_port, QN => n_2904);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n2602, CK => n744, Q => 
                           REGISTERS_29_18_port, QN => n_2905);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n2601, CK => n744, Q => 
                           REGISTERS_29_17_port, QN => n_2906);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n2600, CK => n745, Q => 
                           REGISTERS_29_16_port, QN => n_2907);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n2599, CK => n745, Q => 
                           REGISTERS_29_15_port, QN => n_2908);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n2598, CK => n745, Q => 
                           REGISTERS_29_14_port, QN => n_2909);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n2597, CK => n745, Q => 
                           REGISTERS_29_13_port, QN => n_2910);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n2596, CK => n745, Q => 
                           REGISTERS_29_12_port, QN => n_2911);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n2595, CK => n745, Q => 
                           REGISTERS_29_11_port, QN => n_2912);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n2594, CK => n745, Q => 
                           REGISTERS_29_10_port, QN => n_2913);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n2593, CK => n745, Q => 
                           REGISTERS_29_9_port, QN => n_2914);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n2592, CK => n745, Q => 
                           REGISTERS_29_8_port, QN => n_2915);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n2591, CK => n745, Q => 
                           REGISTERS_29_7_port, QN => n_2916);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n2590, CK => n745, Q => 
                           REGISTERS_29_6_port, QN => n_2917);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n2589, CK => n746, Q => 
                           REGISTERS_29_5_port, QN => n_2918);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n2588, CK => n746, Q => 
                           REGISTERS_29_4_port, QN => n_2919);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n2587, CK => n746, Q => 
                           REGISTERS_29_3_port, QN => n_2920);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n2586, CK => n746, Q => 
                           REGISTERS_29_2_port, QN => n_2921);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n2585, CK => n746, Q => 
                           REGISTERS_29_1_port, QN => n_2922);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n2584, CK => n746, Q => 
                           REGISTERS_29_0_port, QN => n_2923);
   REGISTERS_reg_30_63_inst : DFF_X1 port map( D => n2583, CK => n746, Q => 
                           REGISTERS_30_63_port, QN => n_2924);
   REGISTERS_reg_30_62_inst : DFF_X1 port map( D => n2582, CK => n746, Q => 
                           REGISTERS_30_62_port, QN => n_2925);
   REGISTERS_reg_30_61_inst : DFF_X1 port map( D => n2581, CK => n746, Q => 
                           REGISTERS_30_61_port, QN => n_2926);
   REGISTERS_reg_30_60_inst : DFF_X1 port map( D => n2580, CK => n746, Q => 
                           REGISTERS_30_60_port, QN => n_2927);
   REGISTERS_reg_30_59_inst : DFF_X1 port map( D => n2579, CK => n746, Q => 
                           REGISTERS_30_59_port, QN => n_2928);
   REGISTERS_reg_30_58_inst : DFF_X1 port map( D => n2578, CK => n747, Q => 
                           REGISTERS_30_58_port, QN => n_2929);
   REGISTERS_reg_30_57_inst : DFF_X1 port map( D => n2577, CK => n747, Q => 
                           REGISTERS_30_57_port, QN => n_2930);
   REGISTERS_reg_30_56_inst : DFF_X1 port map( D => n2576, CK => n747, Q => 
                           REGISTERS_30_56_port, QN => n_2931);
   REGISTERS_reg_30_55_inst : DFF_X1 port map( D => n2575, CK => n747, Q => 
                           REGISTERS_30_55_port, QN => n_2932);
   REGISTERS_reg_30_54_inst : DFF_X1 port map( D => n2574, CK => n747, Q => 
                           REGISTERS_30_54_port, QN => n_2933);
   REGISTERS_reg_30_53_inst : DFF_X1 port map( D => n2573, CK => n747, Q => 
                           REGISTERS_30_53_port, QN => n_2934);
   REGISTERS_reg_30_52_inst : DFF_X1 port map( D => n2572, CK => n747, Q => 
                           REGISTERS_30_52_port, QN => n_2935);
   REGISTERS_reg_30_51_inst : DFF_X1 port map( D => n2571, CK => n747, Q => 
                           REGISTERS_30_51_port, QN => n_2936);
   REGISTERS_reg_30_50_inst : DFF_X1 port map( D => n2570, CK => n747, Q => 
                           REGISTERS_30_50_port, QN => n_2937);
   REGISTERS_reg_30_49_inst : DFF_X1 port map( D => n2569, CK => n747, Q => 
                           REGISTERS_30_49_port, QN => n_2938);
   REGISTERS_reg_30_48_inst : DFF_X1 port map( D => n2568, CK => n747, Q => 
                           REGISTERS_30_48_port, QN => n_2939);
   REGISTERS_reg_30_47_inst : DFF_X1 port map( D => n2567, CK => n748, Q => 
                           REGISTERS_30_47_port, QN => n_2940);
   REGISTERS_reg_30_46_inst : DFF_X1 port map( D => n2566, CK => n748, Q => 
                           REGISTERS_30_46_port, QN => n_2941);
   REGISTERS_reg_30_45_inst : DFF_X1 port map( D => n2565, CK => n748, Q => 
                           REGISTERS_30_45_port, QN => n_2942);
   REGISTERS_reg_30_44_inst : DFF_X1 port map( D => n2564, CK => n748, Q => 
                           REGISTERS_30_44_port, QN => n_2943);
   REGISTERS_reg_30_43_inst : DFF_X1 port map( D => n2563, CK => n748, Q => 
                           REGISTERS_30_43_port, QN => n_2944);
   REGISTERS_reg_30_42_inst : DFF_X1 port map( D => n2562, CK => n748, Q => 
                           REGISTERS_30_42_port, QN => n_2945);
   REGISTERS_reg_30_41_inst : DFF_X1 port map( D => n2561, CK => n748, Q => 
                           REGISTERS_30_41_port, QN => n_2946);
   REGISTERS_reg_30_40_inst : DFF_X1 port map( D => n2560, CK => n748, Q => 
                           REGISTERS_30_40_port, QN => n_2947);
   REGISTERS_reg_30_39_inst : DFF_X1 port map( D => n2559, CK => n748, Q => 
                           REGISTERS_30_39_port, QN => n_2948);
   REGISTERS_reg_30_38_inst : DFF_X1 port map( D => n2558, CK => n748, Q => 
                           REGISTERS_30_38_port, QN => n_2949);
   REGISTERS_reg_30_37_inst : DFF_X1 port map( D => n2557, CK => n748, Q => 
                           REGISTERS_30_37_port, QN => n_2950);
   REGISTERS_reg_30_36_inst : DFF_X1 port map( D => n2556, CK => n749, Q => 
                           REGISTERS_30_36_port, QN => n_2951);
   REGISTERS_reg_30_35_inst : DFF_X1 port map( D => n2555, CK => n749, Q => 
                           REGISTERS_30_35_port, QN => n_2952);
   REGISTERS_reg_30_34_inst : DFF_X1 port map( D => n2554, CK => n749, Q => 
                           REGISTERS_30_34_port, QN => n_2953);
   REGISTERS_reg_30_33_inst : DFF_X1 port map( D => n2553, CK => n749, Q => 
                           REGISTERS_30_33_port, QN => n_2954);
   REGISTERS_reg_30_32_inst : DFF_X1 port map( D => n2552, CK => n749, Q => 
                           REGISTERS_30_32_port, QN => n_2955);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n2551, CK => n749, Q => 
                           REGISTERS_30_31_port, QN => n_2956);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n2550, CK => n749, Q => 
                           REGISTERS_30_30_port, QN => n_2957);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n2549, CK => n749, Q => 
                           REGISTERS_30_29_port, QN => n_2958);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n2548, CK => n749, Q => 
                           REGISTERS_30_28_port, QN => n_2959);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n2547, CK => n749, Q => 
                           REGISTERS_30_27_port, QN => n_2960);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n2546, CK => n749, Q => 
                           REGISTERS_30_26_port, QN => n_2961);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n2545, CK => n750, Q => 
                           REGISTERS_30_25_port, QN => n_2962);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n2544, CK => n750, Q => 
                           REGISTERS_30_24_port, QN => n_2963);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n2543, CK => n750, Q => 
                           REGISTERS_30_23_port, QN => n_2964);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n2542, CK => n750, Q => 
                           REGISTERS_30_22_port, QN => n_2965);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n2541, CK => n750, Q => 
                           REGISTERS_30_21_port, QN => n_2966);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n2540, CK => n750, Q => 
                           REGISTERS_30_20_port, QN => n_2967);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n2539, CK => n750, Q => 
                           REGISTERS_30_19_port, QN => n_2968);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n2538, CK => n750, Q => 
                           REGISTERS_30_18_port, QN => n_2969);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n2537, CK => n750, Q => 
                           REGISTERS_30_17_port, QN => n_2970);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n2536, CK => n750, Q => 
                           REGISTERS_30_16_port, QN => n_2971);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n2535, CK => n750, Q => 
                           REGISTERS_30_15_port, QN => n_2972);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n2534, CK => n751, Q => 
                           REGISTERS_30_14_port, QN => n_2973);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n2533, CK => n751, Q => 
                           REGISTERS_30_13_port, QN => n_2974);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n2532, CK => n751, Q => 
                           REGISTERS_30_12_port, QN => n_2975);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n2531, CK => n751, Q => 
                           REGISTERS_30_11_port, QN => n_2976);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n2530, CK => n751, Q => 
                           REGISTERS_30_10_port, QN => n_2977);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n2529, CK => n751, Q => 
                           REGISTERS_30_9_port, QN => n_2978);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n2528, CK => n751, Q => 
                           REGISTERS_30_8_port, QN => n_2979);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n2527, CK => n751, Q => 
                           REGISTERS_30_7_port, QN => n_2980);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n2526, CK => n751, Q => 
                           REGISTERS_30_6_port, QN => n_2981);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n2525, CK => n751, Q => 
                           REGISTERS_30_5_port, QN => n_2982);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n2524, CK => n751, Q => 
                           REGISTERS_30_4_port, QN => n_2983);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n2523, CK => n752, Q => 
                           REGISTERS_30_3_port, QN => n_2984);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n2522, CK => n752, Q => 
                           REGISTERS_30_2_port, QN => n_2985);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n2521, CK => n752, Q => 
                           REGISTERS_30_1_port, QN => n_2986);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n2520, CK => n752, Q => 
                           REGISTERS_30_0_port, QN => n_2987);
   REGISTERS_reg_31_63_inst : DFF_X1 port map( D => n2519, CK => n752, Q => 
                           REGISTERS_31_63_port, QN => n_2988);
   REGISTERS_reg_31_62_inst : DFF_X1 port map( D => n2518, CK => n752, Q => 
                           REGISTERS_31_62_port, QN => n_2989);
   REGISTERS_reg_31_61_inst : DFF_X1 port map( D => n2517, CK => n752, Q => 
                           REGISTERS_31_61_port, QN => n_2990);
   REGISTERS_reg_31_60_inst : DFF_X1 port map( D => n2516, CK => n752, Q => 
                           REGISTERS_31_60_port, QN => n_2991);
   REGISTERS_reg_31_59_inst : DFF_X1 port map( D => n2515, CK => n752, Q => 
                           REGISTERS_31_59_port, QN => n_2992);
   REGISTERS_reg_31_58_inst : DFF_X1 port map( D => n2514, CK => n752, Q => 
                           REGISTERS_31_58_port, QN => n_2993);
   REGISTERS_reg_31_57_inst : DFF_X1 port map( D => n2513, CK => n752, Q => 
                           REGISTERS_31_57_port, QN => n_2994);
   REGISTERS_reg_31_56_inst : DFF_X1 port map( D => n2512, CK => n753, Q => 
                           REGISTERS_31_56_port, QN => n_2995);
   REGISTERS_reg_31_55_inst : DFF_X1 port map( D => n2511, CK => n753, Q => 
                           REGISTERS_31_55_port, QN => n_2996);
   REGISTERS_reg_31_54_inst : DFF_X1 port map( D => n2510, CK => n753, Q => 
                           REGISTERS_31_54_port, QN => n_2997);
   REGISTERS_reg_31_53_inst : DFF_X1 port map( D => n2509, CK => n753, Q => 
                           REGISTERS_31_53_port, QN => n_2998);
   REGISTERS_reg_31_52_inst : DFF_X1 port map( D => n2508, CK => n753, Q => 
                           REGISTERS_31_52_port, QN => n_2999);
   REGISTERS_reg_31_51_inst : DFF_X1 port map( D => n2507, CK => n753, Q => 
                           REGISTERS_31_51_port, QN => n_3000);
   REGISTERS_reg_31_50_inst : DFF_X1 port map( D => n2506, CK => n753, Q => 
                           REGISTERS_31_50_port, QN => n_3001);
   REGISTERS_reg_31_49_inst : DFF_X1 port map( D => n2505, CK => n753, Q => 
                           REGISTERS_31_49_port, QN => n_3002);
   REGISTERS_reg_31_48_inst : DFF_X1 port map( D => n2504, CK => n753, Q => 
                           REGISTERS_31_48_port, QN => n_3003);
   REGISTERS_reg_31_47_inst : DFF_X1 port map( D => n2503, CK => n753, Q => 
                           REGISTERS_31_47_port, QN => n_3004);
   REGISTERS_reg_31_46_inst : DFF_X1 port map( D => n2502, CK => n753, Q => 
                           REGISTERS_31_46_port, QN => n_3005);
   REGISTERS_reg_31_45_inst : DFF_X1 port map( D => n2501, CK => n754, Q => 
                           REGISTERS_31_45_port, QN => n_3006);
   REGISTERS_reg_31_44_inst : DFF_X1 port map( D => n2500, CK => n754, Q => 
                           REGISTERS_31_44_port, QN => n_3007);
   REGISTERS_reg_31_43_inst : DFF_X1 port map( D => n2499, CK => n754, Q => 
                           REGISTERS_31_43_port, QN => n_3008);
   REGISTERS_reg_31_42_inst : DFF_X1 port map( D => n2498, CK => n754, Q => 
                           REGISTERS_31_42_port, QN => n_3009);
   REGISTERS_reg_31_41_inst : DFF_X1 port map( D => n2497, CK => n754, Q => 
                           REGISTERS_31_41_port, QN => n_3010);
   REGISTERS_reg_31_40_inst : DFF_X1 port map( D => n2496, CK => n754, Q => 
                           REGISTERS_31_40_port, QN => n_3011);
   REGISTERS_reg_31_39_inst : DFF_X1 port map( D => n2495, CK => n754, Q => 
                           REGISTERS_31_39_port, QN => n_3012);
   REGISTERS_reg_31_38_inst : DFF_X1 port map( D => n2494, CK => n754, Q => 
                           REGISTERS_31_38_port, QN => n_3013);
   REGISTERS_reg_31_37_inst : DFF_X1 port map( D => n2493, CK => n754, Q => 
                           REGISTERS_31_37_port, QN => n_3014);
   REGISTERS_reg_31_36_inst : DFF_X1 port map( D => n2492, CK => n754, Q => 
                           REGISTERS_31_36_port, QN => n_3015);
   REGISTERS_reg_31_35_inst : DFF_X1 port map( D => n2491, CK => n754, Q => 
                           REGISTERS_31_35_port, QN => n_3016);
   REGISTERS_reg_31_34_inst : DFF_X1 port map( D => n2490, CK => n755, Q => 
                           REGISTERS_31_34_port, QN => n_3017);
   REGISTERS_reg_31_33_inst : DFF_X1 port map( D => n2489, CK => n755, Q => 
                           REGISTERS_31_33_port, QN => n_3018);
   REGISTERS_reg_31_32_inst : DFF_X1 port map( D => n2488, CK => n755, Q => 
                           REGISTERS_31_32_port, QN => n_3019);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n2487, CK => n755, Q => 
                           REGISTERS_31_31_port, QN => n_3020);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n2486, CK => n755, Q => 
                           REGISTERS_31_30_port, QN => n_3021);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n2485, CK => n755, Q => 
                           REGISTERS_31_29_port, QN => n_3022);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n2484, CK => n755, Q => 
                           REGISTERS_31_28_port, QN => n_3023);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n2483, CK => n755, Q => 
                           REGISTERS_31_27_port, QN => n_3024);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n2482, CK => n755, Q => 
                           REGISTERS_31_26_port, QN => n_3025);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n2481, CK => n755, Q => 
                           REGISTERS_31_25_port, QN => n_3026);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n2480, CK => n755, Q => 
                           REGISTERS_31_24_port, QN => n_3027);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n2479, CK => n756, Q => 
                           REGISTERS_31_23_port, QN => n_3028);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n2478, CK => n756, Q => 
                           REGISTERS_31_22_port, QN => n_3029);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n2477, CK => n756, Q => 
                           REGISTERS_31_21_port, QN => n_3030);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n2476, CK => n756, Q => 
                           REGISTERS_31_20_port, QN => n_3031);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n2475, CK => n756, Q => 
                           REGISTERS_31_19_port, QN => n_3032);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n2474, CK => n756, Q => 
                           REGISTERS_31_18_port, QN => n_3033);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n2473, CK => n756, Q => 
                           REGISTERS_31_17_port, QN => n_3034);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n2472, CK => n756, Q => 
                           REGISTERS_31_16_port, QN => n_3035);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n2471, CK => n756, Q => 
                           REGISTERS_31_15_port, QN => n_3036);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n2470, CK => n756, Q => 
                           REGISTERS_31_14_port, QN => n_3037);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n2469, CK => n756, Q => 
                           REGISTERS_31_13_port, QN => n_3038);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n2468, CK => n757, Q => 
                           REGISTERS_31_12_port, QN => n_3039);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n2467, CK => n757, Q => 
                           REGISTERS_31_11_port, QN => n_3040);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n2466, CK => n757, Q => 
                           REGISTERS_31_10_port, QN => n_3041);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n2465, CK => n757, Q => 
                           REGISTERS_31_9_port, QN => n_3042);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n2464, CK => n757, Q => 
                           REGISTERS_31_8_port, QN => n_3043);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n2463, CK => n757, Q => 
                           REGISTERS_31_7_port, QN => n_3044);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n2462, CK => n757, Q => 
                           REGISTERS_31_6_port, QN => n_3045);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n2461, CK => n757, Q => 
                           REGISTERS_31_5_port, QN => n_3046);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n2460, CK => n757, Q => 
                           REGISTERS_31_4_port, QN => n_3047);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n2459, CK => n757, Q => 
                           REGISTERS_31_3_port, QN => n_3048);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n2458, CK => n757, Q => 
                           REGISTERS_31_2_port, QN => n_3049);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n2457, CK => n758, Q => 
                           REGISTERS_31_1_port, QN => n_3050);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n2456, CK => n758, Q => 
                           REGISTERS_31_0_port, QN => n_3051);
   out1_signal_reg_63_inst : DFF_X1 port map( D => n6179, CK => n700, Q => 
                           OUT1(63), QN => n6051);
   out1_signal_reg_62_inst : DFF_X1 port map( D => n6178, CK => n700, Q => 
                           OUT1(62), QN => n6050);
   out1_signal_reg_61_inst : DFF_X1 port map( D => n6177, CK => n700, Q => 
                           OUT1(61), QN => n6049);
   out1_signal_reg_60_inst : DFF_X1 port map( D => n6176, CK => n700, Q => 
                           OUT1(60), QN => n6048);
   out1_signal_reg_59_inst : DFF_X1 port map( D => n6175, CK => n701, Q => 
                           OUT1(59), QN => n6047);
   out1_signal_reg_58_inst : DFF_X1 port map( D => n6174, CK => n701, Q => 
                           OUT1(58), QN => n6046);
   out1_signal_reg_57_inst : DFF_X1 port map( D => n6173, CK => n701, Q => 
                           OUT1(57), QN => n6045);
   out1_signal_reg_56_inst : DFF_X1 port map( D => n6172, CK => n702, Q => 
                           OUT1(56), QN => n6044);
   out1_signal_reg_55_inst : DFF_X1 port map( D => n6171, CK => n702, Q => 
                           OUT1(55), QN => n6043);
   out1_signal_reg_54_inst : DFF_X1 port map( D => n6170, CK => n702, Q => 
                           OUT1(54), QN => n6042);
   out1_signal_reg_53_inst : DFF_X1 port map( D => n6169, CK => n702, Q => 
                           OUT1(53), QN => n6041);
   out1_signal_reg_52_inst : DFF_X1 port map( D => n6168, CK => n703, Q => 
                           OUT1(52), QN => n6040);
   out1_signal_reg_51_inst : DFF_X1 port map( D => n6167, CK => n703, Q => 
                           OUT1(51), QN => n6039);
   out1_signal_reg_50_inst : DFF_X1 port map( D => n6166, CK => n703, Q => 
                           OUT1(50), QN => n6038);
   out1_signal_reg_49_inst : DFF_X1 port map( D => n6165, CK => n703, Q => 
                           OUT1(49), QN => n6037);
   out1_signal_reg_48_inst : DFF_X1 port map( D => n6164, CK => n704, Q => 
                           OUT1(48), QN => n6036);
   out1_signal_reg_47_inst : DFF_X1 port map( D => n6163, CK => n704, Q => 
                           OUT1(47), QN => n6035);
   out1_signal_reg_46_inst : DFF_X1 port map( D => n6162, CK => n704, Q => 
                           OUT1(46), QN => n6034);
   out1_signal_reg_45_inst : DFF_X1 port map( D => n6161, CK => n705, Q => 
                           OUT1(45), QN => n6033);
   out1_signal_reg_44_inst : DFF_X1 port map( D => n6160, CK => n705, Q => 
                           OUT1(44), QN => n6032);
   out1_signal_reg_43_inst : DFF_X1 port map( D => n6159, CK => n705, Q => 
                           OUT1(43), QN => n6031);
   out1_signal_reg_42_inst : DFF_X1 port map( D => n6158, CK => n705, Q => 
                           OUT1(42), QN => n6030);
   out1_signal_reg_41_inst : DFF_X1 port map( D => n6157, CK => n706, Q => 
                           OUT1(41), QN => n6029);
   out1_signal_reg_40_inst : DFF_X1 port map( D => n6156, CK => n706, Q => 
                           OUT1(40), QN => n6028);
   out1_signal_reg_39_inst : DFF_X1 port map( D => n6155, CK => n706, Q => 
                           OUT1(39), QN => n6027);
   out1_signal_reg_38_inst : DFF_X1 port map( D => n6154, CK => n706, Q => 
                           OUT1(38), QN => n6026);
   out1_signal_reg_37_inst : DFF_X1 port map( D => n6153, CK => n707, Q => 
                           OUT1(37), QN => n6025);
   out1_signal_reg_36_inst : DFF_X1 port map( D => n6152, CK => n707, Q => 
                           OUT1(36), QN => n6024);
   out1_signal_reg_35_inst : DFF_X1 port map( D => n6151, CK => n707, Q => 
                           OUT1(35), QN => n6023);
   out1_signal_reg_34_inst : DFF_X1 port map( D => n6150, CK => n708, Q => 
                           OUT1(34), QN => n6022);
   out1_signal_reg_33_inst : DFF_X1 port map( D => n6149, CK => n708, Q => 
                           OUT1(33), QN => n6021);
   out1_signal_reg_32_inst : DFF_X1 port map( D => n6148, CK => n708, Q => 
                           OUT1(32), QN => n6020);
   out1_signal_reg_31_inst : DFF_X1 port map( D => n6147, CK => n708, Q => 
                           OUT1(31), QN => n6019);
   out1_signal_reg_30_inst : DFF_X1 port map( D => n6146, CK => n709, Q => 
                           OUT1(30), QN => n6018);
   out1_signal_reg_29_inst : DFF_X1 port map( D => n6145, CK => n709, Q => 
                           OUT1(29), QN => n6017);
   out1_signal_reg_28_inst : DFF_X1 port map( D => n6144, CK => n709, Q => 
                           OUT1(28), QN => n6016);
   out1_signal_reg_27_inst : DFF_X1 port map( D => n6143, CK => n709, Q => 
                           OUT1(27), QN => n6015);
   out1_signal_reg_26_inst : DFF_X1 port map( D => n6142, CK => n710, Q => 
                           OUT1(26), QN => n6014);
   out1_signal_reg_25_inst : DFF_X1 port map( D => n6141, CK => n710, Q => 
                           OUT1(25), QN => n6013);
   out1_signal_reg_24_inst : DFF_X1 port map( D => n6140, CK => n710, Q => 
                           OUT1(24), QN => n6012);
   out1_signal_reg_23_inst : DFF_X1 port map( D => n6139, CK => n711, Q => 
                           OUT1(23), QN => n6011);
   out1_signal_reg_22_inst : DFF_X1 port map( D => n6138, CK => n711, Q => 
                           OUT1(22), QN => n6010);
   out1_signal_reg_21_inst : DFF_X1 port map( D => n6137, CK => n711, Q => 
                           OUT1(21), QN => n6009);
   out1_signal_reg_20_inst : DFF_X1 port map( D => n6136, CK => n711, Q => 
                           OUT1(20), QN => n6008);
   out1_signal_reg_19_inst : DFF_X1 port map( D => n6135, CK => n712, Q => 
                           OUT1(19), QN => n6007);
   out1_signal_reg_18_inst : DFF_X1 port map( D => n6134, CK => n712, Q => 
                           OUT1(18), QN => n6006);
   out1_signal_reg_17_inst : DFF_X1 port map( D => n6133, CK => n712, Q => 
                           OUT1(17), QN => n6005);
   out1_signal_reg_16_inst : DFF_X1 port map( D => n6132, CK => n712, Q => 
                           OUT1(16), QN => n6004);
   out1_signal_reg_15_inst : DFF_X1 port map( D => n6131, CK => n713, Q => 
                           OUT1(15), QN => n6003);
   out1_signal_reg_14_inst : DFF_X1 port map( D => n6130, CK => n713, Q => 
                           OUT1(14), QN => n6002);
   out1_signal_reg_13_inst : DFF_X1 port map( D => n6129, CK => n713, Q => 
                           OUT1(13), QN => n6001);
   out1_signal_reg_12_inst : DFF_X1 port map( D => n6128, CK => n714, Q => 
                           OUT1(12), QN => n6000);
   out1_signal_reg_11_inst : DFF_X1 port map( D => n6127, CK => n714, Q => 
                           OUT1(11), QN => n5999);
   out1_signal_reg_10_inst : DFF_X1 port map( D => n6126, CK => n714, Q => 
                           OUT1(10), QN => n5998);
   out1_signal_reg_9_inst : DFF_X1 port map( D => n6125, CK => n714, Q => 
                           OUT1(9), QN => n5997);
   out1_signal_reg_8_inst : DFF_X1 port map( D => n6124, CK => n715, Q => 
                           OUT1(8), QN => n5996);
   out1_signal_reg_7_inst : DFF_X1 port map( D => n6123, CK => n715, Q => 
                           OUT1(7), QN => n5995);
   out1_signal_reg_6_inst : DFF_X1 port map( D => n6122, CK => n715, Q => 
                           OUT1(6), QN => n5994);
   out1_signal_reg_5_inst : DFF_X1 port map( D => n6121, CK => n715, Q => 
                           OUT1(5), QN => n5993);
   out1_signal_reg_4_inst : DFF_X1 port map( D => n6120, CK => n716, Q => 
                           OUT1(4), QN => n5992);
   out1_signal_reg_3_inst : DFF_X1 port map( D => n6119, CK => n716, Q => 
                           OUT1(3), QN => n5991);
   out1_signal_reg_2_inst : DFF_X1 port map( D => n6118, CK => n716, Q => 
                           OUT1(2), QN => n5990);
   out1_signal_reg_1_inst : DFF_X1 port map( D => n6117, CK => n717, Q => 
                           OUT1(1), QN => n5989);
   out1_signal_reg_0_inst : DFF_X1 port map( D => n6116, CK => n717, Q => 
                           OUT1(0), QN => n5988);
   out2_signal_reg_63_inst : DFF_X1 port map( D => n6115, CK => n700, Q => 
                           OUT2(63), QN => n5987);
   out2_signal_reg_62_inst : DFF_X1 port map( D => n6114, CK => n700, Q => 
                           OUT2(62), QN => n5986);
   out2_signal_reg_61_inst : DFF_X1 port map( D => n6113, CK => n700, Q => 
                           OUT2(61), QN => n5985);
   out2_signal_reg_60_inst : DFF_X1 port map( D => n6112, CK => n700, Q => 
                           OUT2(60), QN => n5984);
   out2_signal_reg_59_inst : DFF_X1 port map( D => n6111, CK => n701, Q => 
                           OUT2(59), QN => n5983);
   out2_signal_reg_58_inst : DFF_X1 port map( D => n6110, CK => n701, Q => 
                           OUT2(58), QN => n5982);
   out2_signal_reg_57_inst : DFF_X1 port map( D => n6109, CK => n701, Q => 
                           OUT2(57), QN => n5981);
   out2_signal_reg_56_inst : DFF_X1 port map( D => n6108, CK => n701, Q => 
                           OUT2(56), QN => n5980);
   out2_signal_reg_55_inst : DFF_X1 port map( D => n6107, CK => n702, Q => 
                           OUT2(55), QN => n5979);
   out2_signal_reg_54_inst : DFF_X1 port map( D => n6106, CK => n702, Q => 
                           OUT2(54), QN => n5978);
   out2_signal_reg_53_inst : DFF_X1 port map( D => n6105, CK => n702, Q => 
                           OUT2(53), QN => n5977);
   out2_signal_reg_52_inst : DFF_X1 port map( D => n6104, CK => n703, Q => 
                           OUT2(52), QN => n5976);
   out2_signal_reg_51_inst : DFF_X1 port map( D => n6103, CK => n703, Q => 
                           OUT2(51), QN => n5975);
   out2_signal_reg_50_inst : DFF_X1 port map( D => n6102, CK => n703, Q => 
                           OUT2(50), QN => n5974);
   out2_signal_reg_49_inst : DFF_X1 port map( D => n6101, CK => n703, Q => 
                           OUT2(49), QN => n5973);
   out2_signal_reg_48_inst : DFF_X1 port map( D => n6100, CK => n704, Q => 
                           OUT2(48), QN => n5972);
   out2_signal_reg_47_inst : DFF_X1 port map( D => n6099, CK => n704, Q => 
                           OUT2(47), QN => n5971);
   out2_signal_reg_46_inst : DFF_X1 port map( D => n6098, CK => n704, Q => 
                           OUT2(46), QN => n5970);
   out2_signal_reg_45_inst : DFF_X1 port map( D => n6097, CK => n704, Q => 
                           OUT2(45), QN => n5969);
   out2_signal_reg_44_inst : DFF_X1 port map( D => n6096, CK => n705, Q => 
                           OUT2(44), QN => n5968);
   out2_signal_reg_43_inst : DFF_X1 port map( D => n6095, CK => n705, Q => 
                           OUT2(43), QN => n5967);
   out2_signal_reg_42_inst : DFF_X1 port map( D => n6094, CK => n705, Q => 
                           OUT2(42), QN => n5966);
   out2_signal_reg_41_inst : DFF_X1 port map( D => n6093, CK => n706, Q => 
                           OUT2(41), QN => n5965);
   out2_signal_reg_40_inst : DFF_X1 port map( D => n6092, CK => n706, Q => 
                           OUT2(40), QN => n5964);
   out2_signal_reg_39_inst : DFF_X1 port map( D => n6091, CK => n706, Q => 
                           OUT2(39), QN => n5963);
   out2_signal_reg_38_inst : DFF_X1 port map( D => n6090, CK => n706, Q => 
                           OUT2(38), QN => n5962);
   out2_signal_reg_37_inst : DFF_X1 port map( D => n6089, CK => n707, Q => 
                           OUT2(37), QN => n5961);
   out2_signal_reg_36_inst : DFF_X1 port map( D => n6088, CK => n707, Q => 
                           OUT2(36), QN => n5960);
   out2_signal_reg_35_inst : DFF_X1 port map( D => n6087, CK => n707, Q => 
                           OUT2(35), QN => n5959);
   out2_signal_reg_34_inst : DFF_X1 port map( D => n6086, CK => n707, Q => 
                           OUT2(34), QN => n5958);
   out2_signal_reg_33_inst : DFF_X1 port map( D => n6085, CK => n708, Q => 
                           OUT2(33), QN => n5957);
   out2_signal_reg_32_inst : DFF_X1 port map( D => n6084, CK => n708, Q => 
                           OUT2(32), QN => n5956);
   out2_signal_reg_31_inst : DFF_X1 port map( D => n6083, CK => n708, Q => 
                           OUT2(31), QN => n5955);
   out2_signal_reg_30_inst : DFF_X1 port map( D => n6082, CK => n709, Q => 
                           OUT2(30), QN => n5954);
   out2_signal_reg_29_inst : DFF_X1 port map( D => n6081, CK => n709, Q => 
                           OUT2(29), QN => n5953);
   out2_signal_reg_28_inst : DFF_X1 port map( D => n6080, CK => n709, Q => 
                           OUT2(28), QN => n5952);
   out2_signal_reg_27_inst : DFF_X1 port map( D => n6079, CK => n709, Q => 
                           OUT2(27), QN => n5951);
   out2_signal_reg_26_inst : DFF_X1 port map( D => n6078, CK => n710, Q => 
                           OUT2(26), QN => n5950);
   out2_signal_reg_25_inst : DFF_X1 port map( D => n6077, CK => n710, Q => 
                           OUT2(25), QN => n5949);
   out2_signal_reg_24_inst : DFF_X1 port map( D => n6076, CK => n710, Q => 
                           OUT2(24), QN => n5948);
   out2_signal_reg_23_inst : DFF_X1 port map( D => n6075, CK => n710, Q => 
                           OUT2(23), QN => n5947);
   out2_signal_reg_22_inst : DFF_X1 port map( D => n6074, CK => n711, Q => 
                           OUT2(22), QN => n5946);
   out2_signal_reg_21_inst : DFF_X1 port map( D => n6073, CK => n711, Q => 
                           OUT2(21), QN => n5945);
   out2_signal_reg_20_inst : DFF_X1 port map( D => n6072, CK => n711, Q => 
                           OUT2(20), QN => n5944);
   out2_signal_reg_19_inst : DFF_X1 port map( D => n6071, CK => n712, Q => 
                           OUT2(19), QN => n5943);
   out2_signal_reg_18_inst : DFF_X1 port map( D => n6070, CK => n712, Q => 
                           OUT2(18), QN => n5942);
   out2_signal_reg_17_inst : DFF_X1 port map( D => n6069, CK => n712, Q => 
                           OUT2(17), QN => n5941);
   out2_signal_reg_16_inst : DFF_X1 port map( D => n6068, CK => n712, Q => 
                           OUT2(16), QN => n5940);
   out2_signal_reg_15_inst : DFF_X1 port map( D => n6067, CK => n713, Q => 
                           OUT2(15), QN => n5939);
   out2_signal_reg_14_inst : DFF_X1 port map( D => n6066, CK => n713, Q => 
                           OUT2(14), QN => n5938);
   out2_signal_reg_13_inst : DFF_X1 port map( D => n6065, CK => n713, Q => 
                           OUT2(13), QN => n5937);
   out2_signal_reg_12_inst : DFF_X1 port map( D => n6064, CK => n713, Q => 
                           OUT2(12), QN => n5936);
   out2_signal_reg_11_inst : DFF_X1 port map( D => n6063, CK => n714, Q => 
                           OUT2(11), QN => n5935);
   out2_signal_reg_10_inst : DFF_X1 port map( D => n6062, CK => n714, Q => 
                           OUT2(10), QN => n5934);
   out2_signal_reg_9_inst : DFF_X1 port map( D => n6061, CK => n714, Q => 
                           OUT2(9), QN => n5933);
   out2_signal_reg_8_inst : DFF_X1 port map( D => n6060, CK => n715, Q => 
                           OUT2(8), QN => n5932);
   out2_signal_reg_7_inst : DFF_X1 port map( D => n6059, CK => n715, Q => 
                           OUT2(7), QN => n5931);
   out2_signal_reg_6_inst : DFF_X1 port map( D => n6058, CK => n715, Q => 
                           OUT2(6), QN => n5930);
   out2_signal_reg_5_inst : DFF_X1 port map( D => n6057, CK => n715, Q => 
                           OUT2(5), QN => n5929);
   out2_signal_reg_4_inst : DFF_X1 port map( D => n6056, CK => n716, Q => 
                           OUT2(4), QN => n5928);
   out2_signal_reg_3_inst : DFF_X1 port map( D => n6055, CK => n716, Q => 
                           OUT2(3), QN => n5927);
   out2_signal_reg_2_inst : DFF_X1 port map( D => n6054, CK => n716, Q => 
                           OUT2(2), QN => n5926);
   out2_signal_reg_1_inst : DFF_X1 port map( D => n6053, CK => n716, Q => 
                           OUT2(1), QN => n5925);
   out2_signal_reg_0_inst : DFF_X1 port map( D => n6052, CK => n717, Q => 
                           OUT2(0), QN => n5924);
   U3 : OR2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n1);
   U4 : OR2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n2);
   U5 : OR2_X1 port map( A1 => n2276, A2 => ADD_RD1(4), ZN => n3);
   U6 : OR2_X1 port map( A1 => n5678, A2 => ADD_RD2(4), ZN => n4);
   U7 : AND2_X1 port map( A1 => n923, A2 => ADD_RD1(0), ZN => n5);
   U8 : AND2_X1 port map( A1 => n926, A2 => ADD_RD1(0), ZN => n6);
   U9 : AND2_X1 port map( A1 => n925, A2 => ADD_RD1(0), ZN => n7);
   U10 : AND2_X1 port map( A1 => n924, A2 => n2273, ZN => n8);
   U11 : AND2_X1 port map( A1 => n923, A2 => n2273, ZN => n9);
   U12 : AND2_X1 port map( A1 => n926, A2 => n2273, ZN => n10);
   U13 : AND2_X1 port map( A1 => n925, A2 => n2273, ZN => n11);
   U14 : AND2_X1 port map( A1 => n2277, A2 => ADD_RD2(0), ZN => n12);
   U15 : AND2_X1 port map( A1 => n2280, A2 => ADD_RD2(0), ZN => n13);
   U16 : AND2_X1 port map( A1 => n2279, A2 => ADD_RD2(0), ZN => n14);
   U17 : AND2_X1 port map( A1 => n2278, A2 => n5675, ZN => n15);
   U18 : AND2_X1 port map( A1 => n2277, A2 => n5675, ZN => n16);
   U19 : AND2_X1 port map( A1 => n2280, A2 => n5675, ZN => n17);
   U20 : AND2_X1 port map( A1 => n2279, A2 => n5675, ZN => n18);
   U21 : AND2_X1 port map( A1 => ADD_RD1(0), A2 => n924, ZN => n19);
   U22 : AND2_X1 port map( A1 => ADD_RD2(0), A2 => n2278, ZN => n20);
   U23 : OR2_X1 port map( A1 => ENABLE, A2 => RESET, ZN => n21);
   U24 : NAND2_X4 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n5671);
   U25 : AND3_X4 port map( A1 => n692, A2 => n5744, A3 => RD1, ZN => n5746);
   U26 : NAND2_X4 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n2269);
   U27 : NAND2_X4 port map( A1 => ADD_RD2(4), A2 => n5678, ZN => n5673);
   U28 : AND3_X4 port map( A1 => n692, A2 => n5744, A3 => RD2, ZN => n5680);
   U29 : INV_X4 port map( A => n4, ZN => n22);
   U30 : NAND2_X4 port map( A1 => ADD_RD1(4), A2 => n2276, ZN => n2271);
   U31 : INV_X4 port map( A => n2, ZN => n23);
   U32 : INV_X4 port map( A => n3, ZN => n24);
   U33 : INV_X1 port map( A => n5923, ZN => n25);
   U34 : INV_X4 port map( A => n25, ZN => n26);
   U35 : INV_X4 port map( A => n1, ZN => n27);
   U36 : INV_X1 port map( A => n5921, ZN => n28);
   U37 : INV_X4 port map( A => n28, ZN => n29);
   U38 : INV_X1 port map( A => n5922, ZN => n30);
   U39 : INV_X4 port map( A => n30, ZN => n31);
   U40 : INV_X1 port map( A => n5919, ZN => n32);
   U41 : INV_X4 port map( A => n32, ZN => n33);
   U42 : INV_X1 port map( A => n5920, ZN => n34);
   U43 : INV_X4 port map( A => n34, ZN => n35);
   U44 : INV_X1 port map( A => n5917, ZN => n36);
   U45 : INV_X4 port map( A => n36, ZN => n37);
   U46 : INV_X1 port map( A => n5918, ZN => n38);
   U47 : INV_X4 port map( A => n38, ZN => n39);
   U48 : INV_X1 port map( A => n5911, ZN => n40);
   U49 : INV_X4 port map( A => n40, ZN => n41);
   U50 : INV_X1 port map( A => n5912, ZN => n42);
   U51 : INV_X4 port map( A => n42, ZN => n43);
   U52 : INV_X1 port map( A => n5909, ZN => n44);
   U53 : INV_X4 port map( A => n44, ZN => n45);
   U54 : INV_X1 port map( A => n5910, ZN => n46);
   U55 : INV_X4 port map( A => n46, ZN => n47);
   U56 : INV_X1 port map( A => n5907, ZN => n48);
   U57 : INV_X4 port map( A => n48, ZN => n49);
   U58 : INV_X1 port map( A => n5908, ZN => n50);
   U59 : INV_X4 port map( A => n50, ZN => n51);
   U60 : INV_X1 port map( A => n5902, ZN => n52);
   U61 : INV_X4 port map( A => n52, ZN => n53);
   U62 : INV_X1 port map( A => n5903, ZN => n54);
   U63 : INV_X4 port map( A => n54, ZN => n55);
   U64 : INV_X1 port map( A => n5905, ZN => n56);
   U65 : INV_X4 port map( A => n56, ZN => n57);
   U66 : INV_X1 port map( A => n5906, ZN => n58);
   U67 : INV_X4 port map( A => n58, ZN => n59);
   U68 : INV_X1 port map( A => n5898, ZN => n60);
   U69 : INV_X4 port map( A => n60, ZN => n61);
   U70 : INV_X1 port map( A => n5899, ZN => n62);
   U71 : INV_X4 port map( A => n62, ZN => n63);
   U72 : INV_X1 port map( A => n5900, ZN => n64);
   U73 : INV_X4 port map( A => n64, ZN => n65);
   U74 : INV_X1 port map( A => n5901, ZN => n66);
   U75 : INV_X4 port map( A => n66, ZN => n67);
   U76 : INV_X1 port map( A => n5889, ZN => n68);
   U77 : INV_X4 port map( A => n68, ZN => n69);
   U78 : INV_X1 port map( A => n5894, ZN => n70);
   U79 : INV_X4 port map( A => n70, ZN => n71);
   U80 : INV_X1 port map( A => n5896, ZN => n72);
   U81 : INV_X4 port map( A => n72, ZN => n73);
   U82 : INV_X1 port map( A => n5897, ZN => n74);
   U83 : INV_X4 port map( A => n74, ZN => n75);
   U84 : INV_X1 port map( A => n5881, ZN => n76);
   U85 : INV_X4 port map( A => n76, ZN => n77);
   U86 : INV_X1 port map( A => n5883, ZN => n78);
   U87 : INV_X4 port map( A => n78, ZN => n79);
   U88 : INV_X1 port map( A => n5885, ZN => n80);
   U89 : INV_X4 port map( A => n80, ZN => n81);
   U90 : INV_X1 port map( A => n5887, ZN => n82);
   U91 : INV_X4 port map( A => n82, ZN => n83);
   U92 : INV_X1 port map( A => n5811, ZN => n84);
   U93 : INV_X4 port map( A => n84, ZN => n85);
   U94 : INV_X1 port map( A => n5877, ZN => n86);
   U95 : INV_X4 port map( A => n86, ZN => n87);
   U96 : INV_X1 port map( A => n5879, ZN => n88);
   U97 : INV_X4 port map( A => n88, ZN => n89);
   U98 : INV_X4 port map( A => RESET, ZN => n5744);
   U99 : BUF_X1 port map( A => n922, Z => n915);
   U100 : BUF_X1 port map( A => n922, Z => n917);
   U101 : BUF_X1 port map( A => n922, Z => n916);
   U102 : BUF_X1 port map( A => n921, Z => n919);
   U103 : BUF_X1 port map( A => n921, Z => n918);
   U104 : BUF_X1 port map( A => n699, Z => n922);
   U105 : BUF_X1 port map( A => n699, Z => n921);
   U106 : BUF_X1 port map( A => n697, Z => n695);
   U107 : BUF_X1 port map( A => n697, Z => n694);
   U108 : BUF_X1 port map( A => n21, Z => n697);
   U109 : BUF_X1 port map( A => n698, Z => n693);
   U110 : BUF_X1 port map( A => n909, Z => n757);
   U111 : BUF_X1 port map( A => n909, Z => n756);
   U112 : BUF_X1 port map( A => n909, Z => n755);
   U113 : BUF_X1 port map( A => n909, Z => n754);
   U114 : BUF_X1 port map( A => n910, Z => n753);
   U115 : BUF_X1 port map( A => n910, Z => n752);
   U116 : BUF_X1 port map( A => n910, Z => n751);
   U117 : BUF_X1 port map( A => n910, Z => n750);
   U118 : BUF_X1 port map( A => n910, Z => n749);
   U119 : BUF_X1 port map( A => n910, Z => n748);
   U120 : BUF_X1 port map( A => n910, Z => n747);
   U121 : BUF_X1 port map( A => n910, Z => n746);
   U122 : BUF_X1 port map( A => n910, Z => n745);
   U123 : BUF_X1 port map( A => n910, Z => n744);
   U124 : BUF_X1 port map( A => n910, Z => n743);
   U125 : BUF_X1 port map( A => n910, Z => n742);
   U126 : BUF_X1 port map( A => n911, Z => n741);
   U127 : BUF_X1 port map( A => n911, Z => n740);
   U128 : BUF_X1 port map( A => n911, Z => n739);
   U129 : BUF_X1 port map( A => n911, Z => n738);
   U130 : BUF_X1 port map( A => n911, Z => n737);
   U131 : BUF_X1 port map( A => n911, Z => n736);
   U132 : BUF_X1 port map( A => n911, Z => n735);
   U133 : BUF_X1 port map( A => n911, Z => n734);
   U134 : BUF_X1 port map( A => n911, Z => n733);
   U135 : BUF_X1 port map( A => n911, Z => n732);
   U136 : BUF_X1 port map( A => n911, Z => n731);
   U137 : BUF_X1 port map( A => n911, Z => n730);
   U138 : BUF_X1 port map( A => n912, Z => n729);
   U139 : BUF_X1 port map( A => n912, Z => n728);
   U140 : BUF_X1 port map( A => n912, Z => n727);
   U141 : BUF_X1 port map( A => n912, Z => n726);
   U142 : BUF_X1 port map( A => n912, Z => n725);
   U143 : BUF_X1 port map( A => n912, Z => n724);
   U144 : BUF_X1 port map( A => n912, Z => n723);
   U145 : BUF_X1 port map( A => n912, Z => n722);
   U146 : BUF_X1 port map( A => n912, Z => n721);
   U147 : BUF_X1 port map( A => n912, Z => n720);
   U148 : BUF_X1 port map( A => n912, Z => n719);
   U149 : BUF_X1 port map( A => n912, Z => n718);
   U150 : BUF_X1 port map( A => n913, Z => n717);
   U151 : BUF_X1 port map( A => n913, Z => n716);
   U152 : BUF_X1 port map( A => n913, Z => n715);
   U153 : BUF_X1 port map( A => n913, Z => n714);
   U154 : BUF_X1 port map( A => n913, Z => n713);
   U155 : BUF_X1 port map( A => n913, Z => n712);
   U156 : BUF_X1 port map( A => n913, Z => n711);
   U157 : BUF_X1 port map( A => n913, Z => n710);
   U158 : BUF_X1 port map( A => n913, Z => n709);
   U159 : BUF_X1 port map( A => n913, Z => n708);
   U160 : BUF_X1 port map( A => n913, Z => n707);
   U161 : BUF_X1 port map( A => n913, Z => n706);
   U162 : BUF_X1 port map( A => n914, Z => n705);
   U163 : BUF_X1 port map( A => n914, Z => n704);
   U164 : BUF_X1 port map( A => n914, Z => n703);
   U165 : BUF_X1 port map( A => n914, Z => n702);
   U166 : BUF_X1 port map( A => n914, Z => n701);
   U167 : BUF_X1 port map( A => n914, Z => n700);
   U168 : BUF_X1 port map( A => n905, Z => n803);
   U169 : BUF_X1 port map( A => n905, Z => n802);
   U170 : BUF_X1 port map( A => n906, Z => n801);
   U171 : BUF_X1 port map( A => n906, Z => n800);
   U172 : BUF_X1 port map( A => n906, Z => n799);
   U173 : BUF_X1 port map( A => n906, Z => n798);
   U174 : BUF_X1 port map( A => n906, Z => n797);
   U175 : BUF_X1 port map( A => n906, Z => n796);
   U176 : BUF_X1 port map( A => n906, Z => n795);
   U177 : BUF_X1 port map( A => n906, Z => n794);
   U178 : BUF_X1 port map( A => n906, Z => n793);
   U179 : BUF_X1 port map( A => n906, Z => n792);
   U180 : BUF_X1 port map( A => n906, Z => n791);
   U181 : BUF_X1 port map( A => n906, Z => n790);
   U182 : BUF_X1 port map( A => n907, Z => n789);
   U183 : BUF_X1 port map( A => n907, Z => n788);
   U184 : BUF_X1 port map( A => n907, Z => n787);
   U185 : BUF_X1 port map( A => n907, Z => n786);
   U186 : BUF_X1 port map( A => n907, Z => n785);
   U187 : BUF_X1 port map( A => n907, Z => n784);
   U188 : BUF_X1 port map( A => n907, Z => n783);
   U189 : BUF_X1 port map( A => n907, Z => n782);
   U190 : BUF_X1 port map( A => n907, Z => n781);
   U191 : BUF_X1 port map( A => n907, Z => n780);
   U192 : BUF_X1 port map( A => n907, Z => n779);
   U193 : BUF_X1 port map( A => n907, Z => n778);
   U194 : BUF_X1 port map( A => n908, Z => n777);
   U195 : BUF_X1 port map( A => n908, Z => n776);
   U196 : BUF_X1 port map( A => n908, Z => n775);
   U197 : BUF_X1 port map( A => n908, Z => n774);
   U198 : BUF_X1 port map( A => n908, Z => n773);
   U199 : BUF_X1 port map( A => n908, Z => n772);
   U200 : BUF_X1 port map( A => n908, Z => n771);
   U201 : BUF_X1 port map( A => n908, Z => n770);
   U202 : BUF_X1 port map( A => n908, Z => n769);
   U203 : BUF_X1 port map( A => n908, Z => n768);
   U204 : BUF_X1 port map( A => n908, Z => n767);
   U205 : BUF_X1 port map( A => n908, Z => n766);
   U206 : BUF_X1 port map( A => n909, Z => n765);
   U207 : BUF_X1 port map( A => n909, Z => n764);
   U208 : BUF_X1 port map( A => n909, Z => n763);
   U209 : BUF_X1 port map( A => n909, Z => n762);
   U210 : BUF_X1 port map( A => n909, Z => n761);
   U211 : BUF_X1 port map( A => n909, Z => n760);
   U212 : BUF_X1 port map( A => n909, Z => n759);
   U213 : BUF_X1 port map( A => n909, Z => n758);
   U214 : BUF_X1 port map( A => n898, Z => n896);
   U215 : BUF_X1 port map( A => n898, Z => n895);
   U216 : BUF_X1 port map( A => n898, Z => n894);
   U217 : BUF_X1 port map( A => n898, Z => n893);
   U218 : BUF_X1 port map( A => n898, Z => n892);
   U219 : BUF_X1 port map( A => n898, Z => n891);
   U220 : BUF_X1 port map( A => n898, Z => n890);
   U221 : BUF_X1 port map( A => n898, Z => n889);
   U222 : BUF_X1 port map( A => n898, Z => n888);
   U223 : BUF_X1 port map( A => n898, Z => n887);
   U224 : BUF_X1 port map( A => n898, Z => n886);
   U225 : BUF_X1 port map( A => n899, Z => n885);
   U226 : BUF_X1 port map( A => n899, Z => n884);
   U227 : BUF_X1 port map( A => n899, Z => n883);
   U228 : BUF_X1 port map( A => n899, Z => n882);
   U229 : BUF_X1 port map( A => n899, Z => n881);
   U230 : BUF_X1 port map( A => n899, Z => n880);
   U231 : BUF_X1 port map( A => n899, Z => n879);
   U232 : BUF_X1 port map( A => n899, Z => n878);
   U233 : BUF_X1 port map( A => n899, Z => n877);
   U234 : BUF_X1 port map( A => n899, Z => n876);
   U235 : BUF_X1 port map( A => n899, Z => n875);
   U236 : BUF_X1 port map( A => n899, Z => n874);
   U237 : BUF_X1 port map( A => n900, Z => n873);
   U238 : BUF_X1 port map( A => n900, Z => n872);
   U239 : BUF_X1 port map( A => n900, Z => n871);
   U240 : BUF_X1 port map( A => n900, Z => n870);
   U241 : BUF_X1 port map( A => n900, Z => n869);
   U242 : BUF_X1 port map( A => n900, Z => n868);
   U243 : BUF_X1 port map( A => n900, Z => n867);
   U244 : BUF_X1 port map( A => n900, Z => n866);
   U245 : BUF_X1 port map( A => n900, Z => n865);
   U246 : BUF_X1 port map( A => n900, Z => n864);
   U247 : BUF_X1 port map( A => n900, Z => n863);
   U248 : BUF_X1 port map( A => n900, Z => n862);
   U249 : BUF_X1 port map( A => n901, Z => n861);
   U250 : BUF_X1 port map( A => n901, Z => n860);
   U251 : BUF_X1 port map( A => n901, Z => n859);
   U252 : BUF_X1 port map( A => n901, Z => n858);
   U253 : BUF_X1 port map( A => n901, Z => n857);
   U254 : BUF_X1 port map( A => n901, Z => n856);
   U255 : BUF_X1 port map( A => n901, Z => n855);
   U256 : BUF_X1 port map( A => n901, Z => n854);
   U257 : BUF_X1 port map( A => n901, Z => n853);
   U258 : BUF_X1 port map( A => n901, Z => n852);
   U259 : BUF_X1 port map( A => n901, Z => n851);
   U260 : BUF_X1 port map( A => n901, Z => n850);
   U261 : BUF_X1 port map( A => n902, Z => n849);
   U262 : BUF_X1 port map( A => n902, Z => n848);
   U263 : BUF_X1 port map( A => n902, Z => n847);
   U264 : BUF_X1 port map( A => n902, Z => n846);
   U265 : BUF_X1 port map( A => n902, Z => n845);
   U266 : BUF_X1 port map( A => n902, Z => n844);
   U267 : BUF_X1 port map( A => n902, Z => n843);
   U268 : BUF_X1 port map( A => n902, Z => n842);
   U269 : BUF_X1 port map( A => n902, Z => n841);
   U270 : BUF_X1 port map( A => n902, Z => n840);
   U271 : BUF_X1 port map( A => n902, Z => n839);
   U272 : BUF_X1 port map( A => n902, Z => n838);
   U273 : BUF_X1 port map( A => n903, Z => n837);
   U274 : BUF_X1 port map( A => n903, Z => n836);
   U275 : BUF_X1 port map( A => n903, Z => n835);
   U276 : BUF_X1 port map( A => n903, Z => n834);
   U277 : BUF_X1 port map( A => n903, Z => n833);
   U278 : BUF_X1 port map( A => n903, Z => n832);
   U279 : BUF_X1 port map( A => n903, Z => n831);
   U280 : BUF_X1 port map( A => n903, Z => n830);
   U281 : BUF_X1 port map( A => n903, Z => n829);
   U282 : BUF_X1 port map( A => n903, Z => n828);
   U283 : BUF_X1 port map( A => n903, Z => n827);
   U284 : BUF_X1 port map( A => n903, Z => n826);
   U285 : BUF_X1 port map( A => n904, Z => n825);
   U286 : BUF_X1 port map( A => n904, Z => n824);
   U287 : BUF_X1 port map( A => n904, Z => n823);
   U288 : BUF_X1 port map( A => n904, Z => n822);
   U289 : BUF_X1 port map( A => n904, Z => n821);
   U290 : BUF_X1 port map( A => n904, Z => n820);
   U291 : BUF_X1 port map( A => n904, Z => n819);
   U292 : BUF_X1 port map( A => n904, Z => n818);
   U293 : BUF_X1 port map( A => n904, Z => n817);
   U294 : BUF_X1 port map( A => n904, Z => n816);
   U295 : BUF_X1 port map( A => n904, Z => n815);
   U296 : BUF_X1 port map( A => n904, Z => n814);
   U297 : BUF_X1 port map( A => n905, Z => n813);
   U298 : BUF_X1 port map( A => n905, Z => n812);
   U299 : BUF_X1 port map( A => n905, Z => n811);
   U300 : BUF_X1 port map( A => n905, Z => n810);
   U301 : BUF_X1 port map( A => n905, Z => n809);
   U302 : BUF_X1 port map( A => n905, Z => n808);
   U303 : BUF_X1 port map( A => n905, Z => n807);
   U304 : BUF_X1 port map( A => n905, Z => n806);
   U305 : BUF_X1 port map( A => n905, Z => n805);
   U306 : BUF_X1 port map( A => n905, Z => n804);
   U307 : BUF_X1 port map( A => n898, Z => n897);
   U308 : BUF_X1 port map( A => n677, Z => n645);
   U309 : BUF_X1 port map( A => n677, Z => n646);
   U310 : BUF_X1 port map( A => n676, Z => n647);
   U311 : BUF_X1 port map( A => n676, Z => n648);
   U312 : BUF_X1 port map( A => n675, Z => n649);
   U313 : BUF_X1 port map( A => n675, Z => n650);
   U314 : BUF_X1 port map( A => n674, Z => n651);
   U315 : BUF_X1 port map( A => n674, Z => n652);
   U316 : BUF_X1 port map( A => n673, Z => n653);
   U317 : BUF_X1 port map( A => n673, Z => n654);
   U318 : BUF_X1 port map( A => n672, Z => n655);
   U319 : BUF_X1 port map( A => n672, Z => n656);
   U320 : BUF_X1 port map( A => n671, Z => n657);
   U321 : BUF_X1 port map( A => n671, Z => n658);
   U322 : BUF_X1 port map( A => n670, Z => n659);
   U323 : BUF_X1 port map( A => n670, Z => n660);
   U324 : BUF_X1 port map( A => n669, Z => n661);
   U325 : BUF_X1 port map( A => n669, Z => n662);
   U326 : BUF_X1 port map( A => n668, Z => n663);
   U327 : BUF_X1 port map( A => n668, Z => n664);
   U328 : BUF_X1 port map( A => n667, Z => n665);
   U329 : BUF_X1 port map( A => n381, Z => n349);
   U330 : BUF_X1 port map( A => n381, Z => n350);
   U331 : BUF_X1 port map( A => n380, Z => n351);
   U332 : BUF_X1 port map( A => n380, Z => n352);
   U333 : BUF_X1 port map( A => n379, Z => n353);
   U334 : BUF_X1 port map( A => n379, Z => n354);
   U335 : BUF_X1 port map( A => n378, Z => n355);
   U336 : BUF_X1 port map( A => n378, Z => n356);
   U337 : BUF_X1 port map( A => n377, Z => n357);
   U338 : BUF_X1 port map( A => n377, Z => n358);
   U339 : BUF_X1 port map( A => n376, Z => n359);
   U340 : BUF_X1 port map( A => n376, Z => n360);
   U341 : BUF_X1 port map( A => n375, Z => n361);
   U342 : BUF_X1 port map( A => n375, Z => n362);
   U343 : BUF_X1 port map( A => n374, Z => n363);
   U344 : BUF_X1 port map( A => n374, Z => n364);
   U345 : BUF_X1 port map( A => n373, Z => n365);
   U346 : BUF_X1 port map( A => n373, Z => n366);
   U347 : BUF_X1 port map( A => n372, Z => n367);
   U348 : BUF_X1 port map( A => n372, Z => n368);
   U349 : BUF_X1 port map( A => n371, Z => n369);
   U350 : BUF_X1 port map( A => n603, Z => n571);
   U351 : BUF_X1 port map( A => n603, Z => n572);
   U352 : BUF_X1 port map( A => n602, Z => n573);
   U353 : BUF_X1 port map( A => n602, Z => n574);
   U354 : BUF_X1 port map( A => n601, Z => n575);
   U355 : BUF_X1 port map( A => n601, Z => n576);
   U356 : BUF_X1 port map( A => n600, Z => n577);
   U357 : BUF_X1 port map( A => n600, Z => n578);
   U358 : BUF_X1 port map( A => n599, Z => n579);
   U359 : BUF_X1 port map( A => n599, Z => n580);
   U360 : BUF_X1 port map( A => n598, Z => n581);
   U361 : BUF_X1 port map( A => n598, Z => n582);
   U362 : BUF_X1 port map( A => n597, Z => n583);
   U363 : BUF_X1 port map( A => n597, Z => n584);
   U364 : BUF_X1 port map( A => n596, Z => n585);
   U365 : BUF_X1 port map( A => n596, Z => n586);
   U366 : BUF_X1 port map( A => n595, Z => n587);
   U367 : BUF_X1 port map( A => n595, Z => n588);
   U368 : BUF_X1 port map( A => n594, Z => n589);
   U369 : BUF_X1 port map( A => n594, Z => n590);
   U370 : BUF_X1 port map( A => n593, Z => n591);
   U371 : BUF_X1 port map( A => n307, Z => n275_port);
   U372 : BUF_X1 port map( A => n307, Z => n276_port);
   U373 : BUF_X1 port map( A => n306, Z => n277_port);
   U374 : BUF_X1 port map( A => n306, Z => n278_port);
   U375 : BUF_X1 port map( A => n305, Z => n279_port);
   U376 : BUF_X1 port map( A => n305, Z => n280_port);
   U377 : BUF_X1 port map( A => n304, Z => n281_port);
   U378 : BUF_X1 port map( A => n304, Z => n282_port);
   U379 : BUF_X1 port map( A => n303, Z => n283_port);
   U380 : BUF_X1 port map( A => n303, Z => n284_port);
   U381 : BUF_X1 port map( A => n302, Z => n285_port);
   U382 : BUF_X1 port map( A => n302, Z => n286_port);
   U383 : BUF_X1 port map( A => n301, Z => n287_port);
   U384 : BUF_X1 port map( A => n301, Z => n288_port);
   U385 : BUF_X1 port map( A => n300, Z => n289);
   U386 : BUF_X1 port map( A => n300, Z => n290);
   U387 : BUF_X1 port map( A => n299, Z => n291);
   U388 : BUF_X1 port map( A => n299, Z => n292);
   U389 : BUF_X1 port map( A => n298, Z => n293);
   U390 : BUF_X1 port map( A => n298, Z => n294);
   U391 : BUF_X1 port map( A => n297, Z => n295);
   U392 : BUF_X1 port map( A => n640, Z => n608);
   U393 : BUF_X1 port map( A => n640, Z => n609);
   U394 : BUF_X1 port map( A => n639, Z => n610);
   U395 : BUF_X1 port map( A => n639, Z => n611);
   U396 : BUF_X1 port map( A => n638, Z => n612);
   U397 : BUF_X1 port map( A => n638, Z => n613);
   U398 : BUF_X1 port map( A => n637, Z => n614);
   U399 : BUF_X1 port map( A => n637, Z => n615);
   U400 : BUF_X1 port map( A => n636, Z => n616);
   U401 : BUF_X1 port map( A => n636, Z => n617);
   U402 : BUF_X1 port map( A => n635, Z => n618);
   U403 : BUF_X1 port map( A => n635, Z => n619);
   U404 : BUF_X1 port map( A => n634, Z => n620);
   U405 : BUF_X1 port map( A => n634, Z => n621);
   U406 : BUF_X1 port map( A => n633, Z => n622);
   U407 : BUF_X1 port map( A => n633, Z => n623);
   U408 : BUF_X1 port map( A => n632, Z => n624);
   U409 : BUF_X1 port map( A => n632, Z => n625);
   U410 : BUF_X1 port map( A => n631, Z => n626);
   U411 : BUF_X1 port map( A => n631, Z => n627);
   U412 : BUF_X1 port map( A => n630, Z => n628);
   U413 : BUF_X1 port map( A => n344, Z => n312);
   U414 : BUF_X1 port map( A => n344, Z => n313);
   U415 : BUF_X1 port map( A => n343, Z => n314);
   U416 : BUF_X1 port map( A => n343, Z => n315);
   U417 : BUF_X1 port map( A => n342, Z => n316);
   U418 : BUF_X1 port map( A => n342, Z => n317);
   U419 : BUF_X1 port map( A => n341, Z => n318);
   U420 : BUF_X1 port map( A => n341, Z => n319);
   U421 : BUF_X1 port map( A => n340, Z => n320);
   U422 : BUF_X1 port map( A => n340, Z => n321);
   U423 : BUF_X1 port map( A => n339, Z => n322);
   U424 : BUF_X1 port map( A => n339, Z => n323);
   U425 : BUF_X1 port map( A => n338, Z => n324);
   U426 : BUF_X1 port map( A => n338, Z => n325);
   U427 : BUF_X1 port map( A => n337, Z => n326);
   U428 : BUF_X1 port map( A => n337, Z => n327);
   U429 : BUF_X1 port map( A => n336, Z => n328);
   U430 : BUF_X1 port map( A => n336, Z => n329);
   U431 : BUF_X1 port map( A => n335, Z => n330);
   U432 : BUF_X1 port map( A => n335, Z => n331);
   U433 : BUF_X1 port map( A => n334, Z => n332);
   U434 : BUF_X1 port map( A => n566, Z => n534);
   U435 : BUF_X1 port map( A => n566, Z => n535);
   U436 : BUF_X1 port map( A => n565, Z => n536);
   U437 : BUF_X1 port map( A => n565, Z => n537);
   U438 : BUF_X1 port map( A => n564, Z => n538);
   U439 : BUF_X1 port map( A => n564, Z => n539);
   U440 : BUF_X1 port map( A => n563, Z => n540);
   U441 : BUF_X1 port map( A => n563, Z => n541);
   U442 : BUF_X1 port map( A => n562, Z => n542);
   U443 : BUF_X1 port map( A => n562, Z => n543);
   U444 : BUF_X1 port map( A => n561, Z => n544);
   U445 : BUF_X1 port map( A => n561, Z => n545);
   U446 : BUF_X1 port map( A => n560, Z => n546);
   U447 : BUF_X1 port map( A => n560, Z => n547);
   U448 : BUF_X1 port map( A => n559, Z => n548);
   U449 : BUF_X1 port map( A => n559, Z => n549);
   U450 : BUF_X1 port map( A => n558, Z => n550);
   U451 : BUF_X1 port map( A => n558, Z => n551);
   U452 : BUF_X1 port map( A => n557, Z => n552);
   U453 : BUF_X1 port map( A => n557, Z => n553);
   U454 : BUF_X1 port map( A => n556, Z => n554);
   U455 : BUF_X1 port map( A => n270_port, Z => n238_port);
   U456 : BUF_X1 port map( A => n270_port, Z => n239_port);
   U457 : BUF_X1 port map( A => n269_port, Z => n240_port);
   U458 : BUF_X1 port map( A => n269_port, Z => n241_port);
   U459 : BUF_X1 port map( A => n268_port, Z => n242_port);
   U460 : BUF_X1 port map( A => n268_port, Z => n243_port);
   U461 : BUF_X1 port map( A => n267_port, Z => n244_port);
   U462 : BUF_X1 port map( A => n267_port, Z => n245_port);
   U463 : BUF_X1 port map( A => n266_port, Z => n246_port);
   U464 : BUF_X1 port map( A => n266_port, Z => n247_port);
   U465 : BUF_X1 port map( A => n265_port, Z => n248_port);
   U466 : BUF_X1 port map( A => n265_port, Z => n249_port);
   U467 : BUF_X1 port map( A => n264_port, Z => n250_port);
   U468 : BUF_X1 port map( A => n264_port, Z => n251_port);
   U469 : BUF_X1 port map( A => n263_port, Z => n252_port);
   U470 : BUF_X1 port map( A => n263_port, Z => n253_port);
   U471 : BUF_X1 port map( A => n262_port, Z => n254_port);
   U472 : BUF_X1 port map( A => n262_port, Z => n255_port);
   U473 : BUF_X1 port map( A => n261_port, Z => n256_port);
   U474 : BUF_X1 port map( A => n261_port, Z => n257_port);
   U475 : BUF_X1 port map( A => n260_port, Z => n258_port);
   U476 : BUF_X1 port map( A => n916, Z => n910);
   U477 : BUF_X1 port map( A => n916, Z => n911);
   U478 : BUF_X1 port map( A => n915, Z => n912);
   U479 : BUF_X1 port map( A => n915, Z => n913);
   U480 : BUF_X1 port map( A => n917, Z => n906);
   U481 : BUF_X1 port map( A => n917, Z => n907);
   U482 : BUF_X1 port map( A => n917, Z => n908);
   U483 : BUF_X1 port map( A => n916, Z => n909);
   U484 : BUF_X1 port map( A => n919, Z => n900);
   U485 : BUF_X1 port map( A => n919, Z => n901);
   U486 : BUF_X1 port map( A => n919, Z => n902);
   U487 : BUF_X1 port map( A => n918, Z => n903);
   U488 : BUF_X1 port map( A => n918, Z => n904);
   U489 : BUF_X1 port map( A => n918, Z => n905);
   U490 : BUF_X1 port map( A => n920, Z => n898);
   U491 : BUF_X1 port map( A => n920, Z => n899);
   U492 : BUF_X1 port map( A => n915, Z => n914);
   U493 : BUF_X1 port map( A => n667, Z => n666);
   U494 : BUF_X1 port map( A => n371, Z => n370);
   U495 : BUF_X1 port map( A => n593, Z => n592);
   U496 : BUF_X1 port map( A => n297, Z => n296);
   U497 : BUF_X1 port map( A => n630, Z => n629);
   U498 : BUF_X1 port map( A => n334, Z => n333);
   U499 : BUF_X1 port map( A => n556, Z => n555);
   U500 : BUF_X1 port map( A => n260_port, Z => n259_port);
   U501 : BUF_X1 port map( A => n678, Z => n677);
   U502 : BUF_X1 port map( A => n641, Z => n640);
   U503 : BUF_X1 port map( A => n678, Z => n676);
   U504 : BUF_X1 port map( A => n641, Z => n639);
   U505 : BUF_X1 port map( A => n678, Z => n675);
   U506 : BUF_X1 port map( A => n641, Z => n638);
   U507 : BUF_X1 port map( A => n679, Z => n674);
   U508 : BUF_X1 port map( A => n642, Z => n637);
   U509 : BUF_X1 port map( A => n679, Z => n673);
   U510 : BUF_X1 port map( A => n642, Z => n636);
   U511 : BUF_X1 port map( A => n679, Z => n672);
   U512 : BUF_X1 port map( A => n642, Z => n635);
   U513 : BUF_X1 port map( A => n680, Z => n671);
   U514 : BUF_X1 port map( A => n643, Z => n634);
   U515 : BUF_X1 port map( A => n680, Z => n670);
   U516 : BUF_X1 port map( A => n643, Z => n633);
   U517 : BUF_X1 port map( A => n680, Z => n669);
   U518 : BUF_X1 port map( A => n643, Z => n632);
   U519 : BUF_X1 port map( A => n382, Z => n381);
   U520 : BUF_X1 port map( A => n345, Z => n344);
   U521 : BUF_X1 port map( A => n382, Z => n380);
   U522 : BUF_X1 port map( A => n345, Z => n343);
   U523 : BUF_X1 port map( A => n382, Z => n379);
   U524 : BUF_X1 port map( A => n345, Z => n342);
   U525 : BUF_X1 port map( A => n383, Z => n378);
   U526 : BUF_X1 port map( A => n346, Z => n341);
   U527 : BUF_X1 port map( A => n383, Z => n377);
   U528 : BUF_X1 port map( A => n346, Z => n340);
   U529 : BUF_X1 port map( A => n383, Z => n376);
   U530 : BUF_X1 port map( A => n346, Z => n339);
   U531 : BUF_X1 port map( A => n384, Z => n375);
   U532 : BUF_X1 port map( A => n347, Z => n338);
   U533 : BUF_X1 port map( A => n384, Z => n374);
   U534 : BUF_X1 port map( A => n347, Z => n337);
   U535 : BUF_X1 port map( A => n384, Z => n373);
   U536 : BUF_X1 port map( A => n347, Z => n336);
   U537 : BUF_X1 port map( A => n604, Z => n603);
   U538 : BUF_X1 port map( A => n567, Z => n566);
   U539 : BUF_X1 port map( A => n604, Z => n602);
   U540 : BUF_X1 port map( A => n567, Z => n565);
   U541 : BUF_X1 port map( A => n604, Z => n601);
   U542 : BUF_X1 port map( A => n567, Z => n564);
   U543 : BUF_X1 port map( A => n605, Z => n600);
   U544 : BUF_X1 port map( A => n568, Z => n563);
   U545 : BUF_X1 port map( A => n605, Z => n599);
   U546 : BUF_X1 port map( A => n568, Z => n562);
   U547 : BUF_X1 port map( A => n605, Z => n598);
   U548 : BUF_X1 port map( A => n568, Z => n561);
   U549 : BUF_X1 port map( A => n606, Z => n597);
   U550 : BUF_X1 port map( A => n569, Z => n560);
   U551 : BUF_X1 port map( A => n606, Z => n596);
   U552 : BUF_X1 port map( A => n569, Z => n559);
   U553 : BUF_X1 port map( A => n606, Z => n595);
   U554 : BUF_X1 port map( A => n569, Z => n558);
   U555 : BUF_X1 port map( A => n308, Z => n307);
   U556 : BUF_X1 port map( A => n271_port, Z => n270_port);
   U557 : BUF_X1 port map( A => n308, Z => n306);
   U558 : BUF_X1 port map( A => n271_port, Z => n269_port);
   U559 : BUF_X1 port map( A => n308, Z => n305);
   U560 : BUF_X1 port map( A => n271_port, Z => n268_port);
   U561 : BUF_X1 port map( A => n309, Z => n304);
   U562 : BUF_X1 port map( A => n272_port, Z => n267_port);
   U563 : BUF_X1 port map( A => n309, Z => n303);
   U564 : BUF_X1 port map( A => n272_port, Z => n266_port);
   U565 : BUF_X1 port map( A => n309, Z => n302);
   U566 : BUF_X1 port map( A => n272_port, Z => n265_port);
   U567 : BUF_X1 port map( A => n310, Z => n301);
   U568 : BUF_X1 port map( A => n273_port, Z => n264_port);
   U569 : BUF_X1 port map( A => n310, Z => n300);
   U570 : BUF_X1 port map( A => n273_port, Z => n263_port);
   U571 : BUF_X1 port map( A => n310, Z => n299);
   U572 : BUF_X1 port map( A => n273_port, Z => n262_port);
   U573 : BUF_X1 port map( A => n681, Z => n668);
   U574 : BUF_X1 port map( A => n644, Z => n631);
   U575 : BUF_X1 port map( A => n681, Z => n667);
   U576 : BUF_X1 port map( A => n644, Z => n630);
   U577 : BUF_X1 port map( A => n385, Z => n372);
   U578 : BUF_X1 port map( A => n348, Z => n335);
   U579 : BUF_X1 port map( A => n385, Z => n371);
   U580 : BUF_X1 port map( A => n348, Z => n334);
   U581 : BUF_X1 port map( A => n607, Z => n594);
   U582 : BUF_X1 port map( A => n570, Z => n557);
   U583 : BUF_X1 port map( A => n607, Z => n593);
   U584 : BUF_X1 port map( A => n570, Z => n556);
   U585 : BUF_X1 port map( A => n311, Z => n298);
   U586 : BUF_X1 port map( A => n274_port, Z => n261_port);
   U587 : BUF_X1 port map( A => n311, Z => n297);
   U588 : BUF_X1 port map( A => n274_port, Z => n260_port);
   U589 : BUF_X1 port map( A => n921, Z => n920);
   U590 : BUF_X1 port map( A => n529, Z => n497);
   U591 : BUF_X1 port map( A => n455, Z => n423);
   U592 : BUF_X1 port map( A => n529, Z => n498);
   U593 : BUF_X1 port map( A => n455, Z => n424);
   U594 : BUF_X1 port map( A => n528, Z => n499);
   U595 : BUF_X1 port map( A => n454, Z => n425);
   U596 : BUF_X1 port map( A => n528, Z => n500);
   U597 : BUF_X1 port map( A => n454, Z => n426);
   U598 : BUF_X1 port map( A => n527, Z => n501);
   U599 : BUF_X1 port map( A => n453, Z => n427);
   U600 : BUF_X1 port map( A => n527, Z => n502);
   U601 : BUF_X1 port map( A => n453, Z => n428);
   U602 : BUF_X1 port map( A => n526, Z => n503);
   U603 : BUF_X1 port map( A => n452, Z => n429);
   U604 : BUF_X1 port map( A => n526, Z => n504);
   U605 : BUF_X1 port map( A => n452, Z => n430);
   U606 : BUF_X1 port map( A => n525, Z => n505);
   U607 : BUF_X1 port map( A => n451, Z => n431);
   U608 : BUF_X1 port map( A => n525, Z => n506);
   U609 : BUF_X1 port map( A => n451, Z => n432);
   U610 : BUF_X1 port map( A => n524, Z => n507);
   U611 : BUF_X1 port map( A => n450, Z => n433);
   U612 : BUF_X1 port map( A => n524, Z => n508);
   U613 : BUF_X1 port map( A => n450, Z => n434);
   U614 : BUF_X1 port map( A => n523, Z => n509);
   U615 : BUF_X1 port map( A => n449, Z => n435);
   U616 : BUF_X1 port map( A => n523, Z => n510);
   U617 : BUF_X1 port map( A => n449, Z => n436);
   U618 : BUF_X1 port map( A => n522, Z => n511);
   U619 : BUF_X1 port map( A => n448, Z => n437);
   U620 : BUF_X1 port map( A => n522, Z => n512);
   U621 : BUF_X1 port map( A => n448, Z => n438);
   U622 : BUF_X1 port map( A => n521, Z => n513);
   U623 : BUF_X1 port map( A => n447, Z => n439);
   U624 : BUF_X1 port map( A => n521, Z => n514);
   U625 : BUF_X1 port map( A => n447, Z => n440);
   U626 : BUF_X1 port map( A => n520, Z => n515);
   U627 : BUF_X1 port map( A => n446, Z => n441);
   U628 : BUF_X1 port map( A => n520, Z => n516);
   U629 : BUF_X1 port map( A => n446, Z => n442);
   U630 : BUF_X1 port map( A => n519, Z => n517);
   U631 : BUF_X1 port map( A => n445, Z => n443);
   U632 : BUF_X1 port map( A => n233_port, Z => n201);
   U633 : BUF_X1 port map( A => n159_port, Z => n127_port);
   U634 : BUF_X1 port map( A => n233_port, Z => n202);
   U635 : BUF_X1 port map( A => n159_port, Z => n128_port);
   U636 : BUF_X1 port map( A => n232_port, Z => n203);
   U637 : BUF_X1 port map( A => n158_port, Z => n129_port);
   U638 : BUF_X1 port map( A => n232_port, Z => n204);
   U639 : BUF_X1 port map( A => n158_port, Z => n130_port);
   U640 : BUF_X1 port map( A => n231_port, Z => n205);
   U641 : BUF_X1 port map( A => n157_port, Z => n131_port);
   U642 : BUF_X1 port map( A => n231_port, Z => n206);
   U643 : BUF_X1 port map( A => n157_port, Z => n132_port);
   U644 : BUF_X1 port map( A => n230_port, Z => n207);
   U645 : BUF_X1 port map( A => n156_port, Z => n133_port);
   U646 : BUF_X1 port map( A => n230_port, Z => n208);
   U647 : BUF_X1 port map( A => n156_port, Z => n134_port);
   U648 : BUF_X1 port map( A => n229_port, Z => n209);
   U649 : BUF_X1 port map( A => n155_port, Z => n135_port);
   U650 : BUF_X1 port map( A => n229_port, Z => n210);
   U651 : BUF_X1 port map( A => n155_port, Z => n136_port);
   U652 : BUF_X1 port map( A => n228_port, Z => n211);
   U653 : BUF_X1 port map( A => n154_port, Z => n137_port);
   U654 : BUF_X1 port map( A => n228_port, Z => n212);
   U655 : BUF_X1 port map( A => n154_port, Z => n138_port);
   U656 : BUF_X1 port map( A => n227_port, Z => n213);
   U657 : BUF_X1 port map( A => n153_port, Z => n139_port);
   U658 : BUF_X1 port map( A => n227_port, Z => n214);
   U659 : BUF_X1 port map( A => n153_port, Z => n140_port);
   U660 : BUF_X1 port map( A => n226_port, Z => n215);
   U661 : BUF_X1 port map( A => n152_port, Z => n141_port);
   U662 : BUF_X1 port map( A => n226_port, Z => n216);
   U663 : BUF_X1 port map( A => n152_port, Z => n142_port);
   U664 : BUF_X1 port map( A => n225_port, Z => n217);
   U665 : BUF_X1 port map( A => n151_port, Z => n143_port);
   U666 : BUF_X1 port map( A => n225_port, Z => n218);
   U667 : BUF_X1 port map( A => n151_port, Z => n144_port);
   U668 : BUF_X1 port map( A => n224, Z => n219);
   U669 : BUF_X1 port map( A => n150_port, Z => n145_port);
   U670 : BUF_X1 port map( A => n224, Z => n220);
   U671 : BUF_X1 port map( A => n150_port, Z => n146_port);
   U672 : BUF_X1 port map( A => n223, Z => n221);
   U673 : BUF_X1 port map( A => n149_port, Z => n147_port);
   U674 : BUF_X1 port map( A => n492, Z => n460);
   U675 : BUF_X1 port map( A => n418, Z => n386);
   U676 : BUF_X1 port map( A => n492, Z => n461);
   U677 : BUF_X1 port map( A => n418, Z => n387);
   U678 : BUF_X1 port map( A => n491, Z => n462);
   U679 : BUF_X1 port map( A => n417, Z => n388);
   U680 : BUF_X1 port map( A => n491, Z => n463);
   U681 : BUF_X1 port map( A => n417, Z => n389);
   U682 : BUF_X1 port map( A => n490, Z => n464);
   U683 : BUF_X1 port map( A => n416, Z => n390);
   U684 : BUF_X1 port map( A => n490, Z => n465);
   U685 : BUF_X1 port map( A => n416, Z => n391);
   U686 : BUF_X1 port map( A => n489, Z => n466);
   U687 : BUF_X1 port map( A => n415, Z => n392);
   U688 : BUF_X1 port map( A => n489, Z => n467);
   U689 : BUF_X1 port map( A => n415, Z => n393);
   U690 : BUF_X1 port map( A => n488, Z => n468);
   U691 : BUF_X1 port map( A => n414, Z => n394);
   U692 : BUF_X1 port map( A => n488, Z => n469);
   U693 : BUF_X1 port map( A => n414, Z => n395);
   U694 : BUF_X1 port map( A => n487, Z => n470);
   U695 : BUF_X1 port map( A => n413, Z => n396);
   U696 : BUF_X1 port map( A => n487, Z => n471);
   U697 : BUF_X1 port map( A => n413, Z => n397);
   U698 : BUF_X1 port map( A => n486, Z => n472);
   U699 : BUF_X1 port map( A => n412, Z => n398);
   U700 : BUF_X1 port map( A => n486, Z => n473);
   U701 : BUF_X1 port map( A => n412, Z => n399);
   U702 : BUF_X1 port map( A => n485, Z => n474);
   U703 : BUF_X1 port map( A => n411, Z => n400);
   U704 : BUF_X1 port map( A => n485, Z => n475);
   U705 : BUF_X1 port map( A => n411, Z => n401);
   U706 : BUF_X1 port map( A => n484, Z => n476);
   U707 : BUF_X1 port map( A => n410, Z => n402);
   U708 : BUF_X1 port map( A => n484, Z => n477);
   U709 : BUF_X1 port map( A => n410, Z => n403);
   U710 : BUF_X1 port map( A => n483, Z => n478);
   U711 : BUF_X1 port map( A => n409, Z => n404);
   U712 : BUF_X1 port map( A => n483, Z => n479);
   U713 : BUF_X1 port map( A => n409, Z => n405);
   U714 : BUF_X1 port map( A => n482, Z => n480);
   U715 : BUF_X1 port map( A => n408, Z => n406);
   U716 : BUF_X1 port map( A => n196, Z => n164);
   U717 : BUF_X1 port map( A => n122_port, Z => n90);
   U718 : BUF_X1 port map( A => n196, Z => n165);
   U719 : BUF_X1 port map( A => n122_port, Z => n91);
   U720 : BUF_X1 port map( A => n195, Z => n166);
   U721 : BUF_X1 port map( A => n121_port, Z => n92);
   U722 : BUF_X1 port map( A => n195, Z => n167);
   U723 : BUF_X1 port map( A => n121_port, Z => n93);
   U724 : BUF_X1 port map( A => n194, Z => n168);
   U725 : BUF_X1 port map( A => n120_port, Z => n94);
   U726 : BUF_X1 port map( A => n194, Z => n169);
   U727 : BUF_X1 port map( A => n120_port, Z => n95);
   U728 : BUF_X1 port map( A => n193, Z => n170);
   U729 : BUF_X1 port map( A => n119_port, Z => n96_port);
   U730 : BUF_X1 port map( A => n193, Z => n171);
   U731 : BUF_X1 port map( A => n119_port, Z => n97_port);
   U732 : BUF_X1 port map( A => n192, Z => n172);
   U733 : BUF_X1 port map( A => n118_port, Z => n98_port);
   U734 : BUF_X1 port map( A => n192, Z => n173);
   U735 : BUF_X1 port map( A => n118_port, Z => n99_port);
   U736 : BUF_X1 port map( A => n191, Z => n174);
   U737 : BUF_X1 port map( A => n117_port, Z => n100_port);
   U738 : BUF_X1 port map( A => n191, Z => n175);
   U739 : BUF_X1 port map( A => n117_port, Z => n101_port);
   U740 : BUF_X1 port map( A => n190, Z => n176);
   U741 : BUF_X1 port map( A => n116_port, Z => n102_port);
   U742 : BUF_X1 port map( A => n190, Z => n177);
   U743 : BUF_X1 port map( A => n116_port, Z => n103_port);
   U744 : BUF_X1 port map( A => n189, Z => n178);
   U745 : BUF_X1 port map( A => n115_port, Z => n104_port);
   U746 : BUF_X1 port map( A => n189, Z => n179);
   U747 : BUF_X1 port map( A => n115_port, Z => n105_port);
   U748 : BUF_X1 port map( A => n188, Z => n180);
   U749 : BUF_X1 port map( A => n114_port, Z => n106_port);
   U750 : BUF_X1 port map( A => n188, Z => n181);
   U751 : BUF_X1 port map( A => n114_port, Z => n107_port);
   U752 : BUF_X1 port map( A => n187, Z => n182);
   U753 : BUF_X1 port map( A => n113_port, Z => n108_port);
   U754 : BUF_X1 port map( A => n187, Z => n183);
   U755 : BUF_X1 port map( A => n113_port, Z => n109_port);
   U756 : BUF_X1 port map( A => n186, Z => n184);
   U757 : BUF_X1 port map( A => n112_port, Z => n110_port);
   U758 : BUF_X1 port map( A => n695, Z => n684);
   U759 : BUF_X1 port map( A => n695, Z => n685);
   U760 : BUF_X1 port map( A => n695, Z => n686);
   U761 : BUF_X1 port map( A => n694, Z => n687);
   U762 : BUF_X1 port map( A => n694, Z => n688);
   U763 : BUF_X1 port map( A => n694, Z => n689);
   U764 : BUF_X1 port map( A => n696, Z => n682);
   U765 : BUF_X1 port map( A => n696, Z => n683);
   U766 : BUF_X1 port map( A => n519, Z => n518);
   U767 : BUF_X1 port map( A => n445, Z => n444);
   U768 : BUF_X1 port map( A => n223, Z => n222);
   U769 : BUF_X1 port map( A => n149_port, Z => n148_port);
   U770 : BUF_X1 port map( A => n482, Z => n481);
   U771 : BUF_X1 port map( A => n408, Z => n407);
   U772 : BUF_X1 port map( A => n186, Z => n185);
   U773 : BUF_X1 port map( A => n112_port, Z => n111_port);
   U774 : BUF_X1 port map( A => n530, Z => n529);
   U775 : BUF_X1 port map( A => n493, Z => n492);
   U776 : BUF_X1 port map( A => n456, Z => n455);
   U777 : BUF_X1 port map( A => n419, Z => n418);
   U778 : BUF_X1 port map( A => n530, Z => n528);
   U779 : BUF_X1 port map( A => n493, Z => n491);
   U780 : BUF_X1 port map( A => n456, Z => n454);
   U781 : BUF_X1 port map( A => n419, Z => n417);
   U782 : BUF_X1 port map( A => n530, Z => n527);
   U783 : BUF_X1 port map( A => n493, Z => n490);
   U784 : BUF_X1 port map( A => n456, Z => n453);
   U785 : BUF_X1 port map( A => n419, Z => n416);
   U786 : BUF_X1 port map( A => n531, Z => n526);
   U787 : BUF_X1 port map( A => n494, Z => n489);
   U788 : BUF_X1 port map( A => n457, Z => n452);
   U789 : BUF_X1 port map( A => n420, Z => n415);
   U790 : BUF_X1 port map( A => n531, Z => n525);
   U791 : BUF_X1 port map( A => n494, Z => n488);
   U792 : BUF_X1 port map( A => n457, Z => n451);
   U793 : BUF_X1 port map( A => n420, Z => n414);
   U794 : BUF_X1 port map( A => n531, Z => n524);
   U795 : BUF_X1 port map( A => n494, Z => n487);
   U796 : BUF_X1 port map( A => n457, Z => n450);
   U797 : BUF_X1 port map( A => n420, Z => n413);
   U798 : BUF_X1 port map( A => n532, Z => n523);
   U799 : BUF_X1 port map( A => n495, Z => n486);
   U800 : BUF_X1 port map( A => n458, Z => n449);
   U801 : BUF_X1 port map( A => n421, Z => n412);
   U802 : BUF_X1 port map( A => n532, Z => n522);
   U803 : BUF_X1 port map( A => n495, Z => n485);
   U804 : BUF_X1 port map( A => n458, Z => n448);
   U805 : BUF_X1 port map( A => n421, Z => n411);
   U806 : BUF_X1 port map( A => n532, Z => n521);
   U807 : BUF_X1 port map( A => n495, Z => n484);
   U808 : BUF_X1 port map( A => n458, Z => n447);
   U809 : BUF_X1 port map( A => n421, Z => n410);
   U810 : BUF_X1 port map( A => n234_port, Z => n233_port);
   U811 : BUF_X1 port map( A => n197, Z => n196);
   U812 : BUF_X1 port map( A => n160, Z => n159_port);
   U813 : BUF_X1 port map( A => n123_port, Z => n122_port);
   U814 : BUF_X1 port map( A => n234_port, Z => n232_port);
   U815 : BUF_X1 port map( A => n197, Z => n195);
   U816 : BUF_X1 port map( A => n160, Z => n158_port);
   U817 : BUF_X1 port map( A => n123_port, Z => n121_port);
   U818 : BUF_X1 port map( A => n234_port, Z => n231_port);
   U819 : BUF_X1 port map( A => n197, Z => n194);
   U820 : BUF_X1 port map( A => n160, Z => n157_port);
   U821 : BUF_X1 port map( A => n123_port, Z => n120_port);
   U822 : BUF_X1 port map( A => n235_port, Z => n230_port);
   U823 : BUF_X1 port map( A => n198, Z => n193);
   U824 : BUF_X1 port map( A => n161, Z => n156_port);
   U825 : BUF_X1 port map( A => n124_port, Z => n119_port);
   U826 : BUF_X1 port map( A => n235_port, Z => n229_port);
   U827 : BUF_X1 port map( A => n198, Z => n192);
   U828 : BUF_X1 port map( A => n161, Z => n155_port);
   U829 : BUF_X1 port map( A => n124_port, Z => n118_port);
   U830 : BUF_X1 port map( A => n235_port, Z => n228_port);
   U831 : BUF_X1 port map( A => n198, Z => n191);
   U832 : BUF_X1 port map( A => n161, Z => n154_port);
   U833 : BUF_X1 port map( A => n124_port, Z => n117_port);
   U834 : BUF_X1 port map( A => n236_port, Z => n227_port);
   U835 : BUF_X1 port map( A => n199, Z => n190);
   U836 : BUF_X1 port map( A => n162, Z => n153_port);
   U837 : BUF_X1 port map( A => n125_port, Z => n116_port);
   U838 : BUF_X1 port map( A => n236_port, Z => n226_port);
   U839 : BUF_X1 port map( A => n199, Z => n189);
   U840 : BUF_X1 port map( A => n162, Z => n152_port);
   U841 : BUF_X1 port map( A => n125_port, Z => n115_port);
   U842 : BUF_X1 port map( A => n236_port, Z => n225_port);
   U843 : BUF_X1 port map( A => n199, Z => n188);
   U844 : BUF_X1 port map( A => n162, Z => n151_port);
   U845 : BUF_X1 port map( A => n125_port, Z => n114_port);
   U846 : BUF_X1 port map( A => n533, Z => n520);
   U847 : BUF_X1 port map( A => n496, Z => n483);
   U848 : BUF_X1 port map( A => n459, Z => n446);
   U849 : BUF_X1 port map( A => n422, Z => n409);
   U850 : BUF_X1 port map( A => n533, Z => n519);
   U851 : BUF_X1 port map( A => n496, Z => n482);
   U852 : BUF_X1 port map( A => n459, Z => n445);
   U853 : BUF_X1 port map( A => n422, Z => n408);
   U854 : BUF_X1 port map( A => n237_port, Z => n224);
   U855 : BUF_X1 port map( A => n200, Z => n187);
   U856 : BUF_X1 port map( A => n163, Z => n150_port);
   U857 : BUF_X1 port map( A => n126_port, Z => n113_port);
   U858 : BUF_X1 port map( A => n237_port, Z => n223);
   U859 : BUF_X1 port map( A => n200, Z => n186);
   U860 : BUF_X1 port map( A => n163, Z => n149_port);
   U861 : BUF_X1 port map( A => n126_port, Z => n112_port);
   U862 : BUF_X1 port map( A => n18, Z => n678);
   U863 : BUF_X1 port map( A => n17, Z => n641);
   U864 : BUF_X1 port map( A => n18, Z => n679);
   U865 : BUF_X1 port map( A => n17, Z => n642);
   U866 : BUF_X1 port map( A => n18, Z => n680);
   U867 : BUF_X1 port map( A => n17, Z => n643);
   U868 : BUF_X1 port map( A => n11, Z => n382);
   U869 : BUF_X1 port map( A => n10, Z => n345);
   U870 : BUF_X1 port map( A => n11, Z => n383);
   U871 : BUF_X1 port map( A => n10, Z => n346);
   U872 : BUF_X1 port map( A => n11, Z => n384);
   U873 : BUF_X1 port map( A => n10, Z => n347);
   U874 : BUF_X1 port map( A => n16, Z => n604);
   U875 : BUF_X1 port map( A => n15, Z => n567);
   U876 : BUF_X1 port map( A => n16, Z => n605);
   U877 : BUF_X1 port map( A => n15, Z => n568);
   U878 : BUF_X1 port map( A => n16, Z => n606);
   U879 : BUF_X1 port map( A => n15, Z => n569);
   U880 : BUF_X1 port map( A => n9, Z => n308);
   U881 : BUF_X1 port map( A => n8, Z => n271_port);
   U882 : BUF_X1 port map( A => n9, Z => n309);
   U883 : BUF_X1 port map( A => n8, Z => n272_port);
   U884 : BUF_X1 port map( A => n9, Z => n310);
   U885 : BUF_X1 port map( A => n8, Z => n273_port);
   U886 : BUF_X1 port map( A => n697, Z => n696);
   U887 : BUF_X1 port map( A => n18, Z => n681);
   U888 : BUF_X1 port map( A => n17, Z => n644);
   U889 : BUF_X1 port map( A => n11, Z => n385);
   U890 : BUF_X1 port map( A => n10, Z => n348);
   U891 : BUF_X1 port map( A => n16, Z => n607);
   U892 : BUF_X1 port map( A => n15, Z => n570);
   U893 : BUF_X1 port map( A => n9, Z => n311);
   U894 : BUF_X1 port map( A => n8, Z => n274_port);
   U895 : BUF_X1 port map( A => n693, Z => n690);
   U896 : BUF_X1 port map( A => n693, Z => n691);
   U897 : BUF_X1 port map( A => n693, Z => n692);
   U898 : INV_X1 port map( A => ADD_RD2(1), ZN => n5676);
   U899 : INV_X1 port map( A => ADD_RD1(1), ZN => n2274);
   U900 : INV_X1 port map( A => ADD_RD2(3), ZN => n5678);
   U901 : INV_X1 port map( A => ADD_RD1(3), ZN => n2276);
   U902 : INV_X1 port map( A => ADD_RD2(2), ZN => n5677);
   U903 : INV_X1 port map( A => ADD_RD1(2), ZN => n2275);
   U904 : BUF_X1 port map( A => n21, Z => n698);
   U905 : BUF_X1 port map( A => n14, Z => n530);
   U906 : BUF_X1 port map( A => n13, Z => n493);
   U907 : BUF_X1 port map( A => n12, Z => n456);
   U908 : BUF_X1 port map( A => n20, Z => n419);
   U909 : BUF_X1 port map( A => n14, Z => n531);
   U910 : BUF_X1 port map( A => n13, Z => n494);
   U911 : BUF_X1 port map( A => n12, Z => n457);
   U912 : BUF_X1 port map( A => n20, Z => n420);
   U913 : BUF_X1 port map( A => n14, Z => n532);
   U914 : BUF_X1 port map( A => n13, Z => n495);
   U915 : BUF_X1 port map( A => n12, Z => n458);
   U916 : BUF_X1 port map( A => n20, Z => n421);
   U917 : BUF_X1 port map( A => n7, Z => n234_port);
   U918 : BUF_X1 port map( A => n6, Z => n197);
   U919 : BUF_X1 port map( A => n5, Z => n160);
   U920 : BUF_X1 port map( A => n19, Z => n123_port);
   U921 : BUF_X1 port map( A => n7, Z => n235_port);
   U922 : BUF_X1 port map( A => n6, Z => n198);
   U923 : BUF_X1 port map( A => n5, Z => n161);
   U924 : BUF_X1 port map( A => n19, Z => n124_port);
   U925 : BUF_X1 port map( A => n7, Z => n236_port);
   U926 : BUF_X1 port map( A => n6, Z => n199);
   U927 : BUF_X1 port map( A => n5, Z => n162);
   U928 : BUF_X1 port map( A => n19, Z => n125_port);
   U929 : BUF_X1 port map( A => CLK, Z => n699);
   U930 : BUF_X1 port map( A => n14, Z => n533);
   U931 : BUF_X1 port map( A => n13, Z => n496);
   U932 : BUF_X1 port map( A => n12, Z => n459);
   U933 : BUF_X1 port map( A => n20, Z => n422);
   U934 : BUF_X1 port map( A => n7, Z => n237_port);
   U935 : BUF_X1 port map( A => n6, Z => n200);
   U936 : BUF_X1 port map( A => n5, Z => n163);
   U937 : BUF_X1 port map( A => n19, Z => n126_port);
   U938 : INV_X1 port map( A => ADD_RD2(0), ZN => n5675);
   U939 : INV_X1 port map( A => ADD_RD1(0), ZN => n2273);
   U940 : NOR2_X1 port map( A1 => n2275, A2 => ADD_RD1(1), ZN => n923);
   U941 : NOR2_X1 port map( A1 => n2275, A2 => n2274, ZN => n924);
   U942 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n127_port, B1 => 
                           REGISTERS_23_0_port, B2 => n90, ZN => n930);
   U943 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n925);
   U944 : NOR2_X1 port map( A1 => n2274, A2 => ADD_RD1(2), ZN => n926);
   U945 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n201, B1 => 
                           REGISTERS_19_0_port, B2 => n164, ZN => n929);
   U946 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n275_port, B1 => 
                           REGISTERS_22_0_port, B2 => n238_port, ZN => n928);
   U947 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n349, B1 => 
                           REGISTERS_18_0_port, B2 => n312, ZN => n927);
   U948 : AND4_X1 port map( A1 => n930, A2 => n929, A3 => n928, A4 => n927, ZN 
                           => n947);
   U949 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n127_port, B1 => 
                           REGISTERS_31_0_port, B2 => n90, ZN => n934);
   U950 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n201, B1 => 
                           REGISTERS_27_0_port, B2 => n164, ZN => n933);
   U951 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n275_port, B1 => 
                           REGISTERS_30_0_port, B2 => n238_port, ZN => n932);
   U952 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n349, B1 => 
                           REGISTERS_26_0_port, B2 => n312, ZN => n931);
   U953 : AND4_X1 port map( A1 => n934, A2 => n933, A3 => n932, A4 => n931, ZN 
                           => n946);
   U954 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n127_port, B1 => 
                           REGISTERS_7_0_port, B2 => n90, ZN => n938);
   U955 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n201, B1 => 
                           REGISTERS_3_0_port, B2 => n164, ZN => n937);
   U956 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n275_port, B1 => 
                           REGISTERS_6_0_port, B2 => n238_port, ZN => n936);
   U957 : AOI22_X1 port map( A1 => REGISTERS_0_0_port, A2 => n349, B1 => 
                           REGISTERS_2_0_port, B2 => n312, ZN => n935);
   U958 : NAND4_X1 port map( A1 => n938, A2 => n937, A3 => n936, A4 => n935, ZN
                           => n944);
   U959 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n127_port, B1 => 
                           REGISTERS_15_0_port, B2 => n90, ZN => n942);
   U960 : AOI22_X1 port map( A1 => REGISTERS_9_0_port, A2 => n201, B1 => 
                           REGISTERS_11_0_port, B2 => n164, ZN => n941);
   U961 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n275_port, B1 => 
                           REGISTERS_14_0_port, B2 => n238_port, ZN => n940);
   U962 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n349, B1 => 
                           REGISTERS_10_0_port, B2 => n312, ZN => n939);
   U963 : NAND4_X1 port map( A1 => n942, A2 => n941, A3 => n940, A4 => n939, ZN
                           => n943);
   U964 : AOI22_X1 port map( A1 => n944, A2 => n27, B1 => n943, B2 => n24, ZN 
                           => n945);
   U965 : OAI221_X1 port map( B1 => n2271, B2 => n947, C1 => n2269, C2 => n946,
                           A => n945, ZN => N159);
   U966 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n127_port, B1 => 
                           REGISTERS_23_1_port, B2 => n90, ZN => n951);
   U967 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n201, B1 => 
                           REGISTERS_19_1_port, B2 => n164, ZN => n950);
   U968 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n275_port, B1 => 
                           REGISTERS_22_1_port, B2 => n238_port, ZN => n949);
   U969 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n349, B1 => 
                           REGISTERS_18_1_port, B2 => n312, ZN => n948);
   U970 : AND4_X1 port map( A1 => n951, A2 => n950, A3 => n949, A4 => n948, ZN 
                           => n968);
   U971 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n127_port, B1 => 
                           REGISTERS_31_1_port, B2 => n90, ZN => n955);
   U972 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n201, B1 => 
                           REGISTERS_27_1_port, B2 => n164, ZN => n954);
   U973 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n275_port, B1 => 
                           REGISTERS_30_1_port, B2 => n238_port, ZN => n953);
   U974 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n349, B1 => 
                           REGISTERS_26_1_port, B2 => n312, ZN => n952);
   U975 : AND4_X1 port map( A1 => n955, A2 => n954, A3 => n953, A4 => n952, ZN 
                           => n967);
   U976 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n127_port, B1 => 
                           REGISTERS_7_1_port, B2 => n90, ZN => n959);
   U977 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n201, B1 => 
                           REGISTERS_3_1_port, B2 => n164, ZN => n958);
   U978 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n275_port, B1 => 
                           REGISTERS_6_1_port, B2 => n238_port, ZN => n957);
   U979 : AOI22_X1 port map( A1 => REGISTERS_0_1_port, A2 => n349, B1 => 
                           REGISTERS_2_1_port, B2 => n312, ZN => n956);
   U980 : NAND4_X1 port map( A1 => n959, A2 => n958, A3 => n957, A4 => n956, ZN
                           => n965);
   U981 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n127_port, B1 => 
                           REGISTERS_15_1_port, B2 => n90, ZN => n963);
   U982 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n201, B1 => 
                           REGISTERS_11_1_port, B2 => n164, ZN => n962);
   U983 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n275_port, B1 => 
                           REGISTERS_14_1_port, B2 => n238_port, ZN => n961);
   U984 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n349, B1 => 
                           REGISTERS_10_1_port, B2 => n312, ZN => n960);
   U985 : NAND4_X1 port map( A1 => n963, A2 => n962, A3 => n961, A4 => n960, ZN
                           => n964);
   U986 : AOI22_X1 port map( A1 => n965, A2 => n27, B1 => n964, B2 => n24, ZN 
                           => n966);
   U987 : OAI221_X1 port map( B1 => n2271, B2 => n968, C1 => n2269, C2 => n967,
                           A => n966, ZN => N158);
   U988 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n127_port, B1 => 
                           REGISTERS_23_2_port, B2 => n90, ZN => n972);
   U989 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n201, B1 => 
                           REGISTERS_19_2_port, B2 => n164, ZN => n971);
   U990 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n275_port, B1 => 
                           REGISTERS_22_2_port, B2 => n238_port, ZN => n970);
   U991 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n349, B1 => 
                           REGISTERS_18_2_port, B2 => n312, ZN => n969);
   U992 : AND4_X1 port map( A1 => n972, A2 => n971, A3 => n970, A4 => n969, ZN 
                           => n989);
   U993 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n127_port, B1 => 
                           REGISTERS_31_2_port, B2 => n90, ZN => n976);
   U994 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n201, B1 => 
                           REGISTERS_27_2_port, B2 => n164, ZN => n975);
   U995 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n275_port, B1 => 
                           REGISTERS_30_2_port, B2 => n238_port, ZN => n974);
   U996 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n349, B1 => 
                           REGISTERS_26_2_port, B2 => n312, ZN => n973);
   U997 : AND4_X1 port map( A1 => n976, A2 => n975, A3 => n974, A4 => n973, ZN 
                           => n988);
   U998 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n127_port, B1 => 
                           REGISTERS_7_2_port, B2 => n90, ZN => n980);
   U999 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n201, B1 => 
                           REGISTERS_3_2_port, B2 => n164, ZN => n979);
   U1000 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n275_port, B1 => 
                           REGISTERS_6_2_port, B2 => n238_port, ZN => n978);
   U1001 : AOI22_X1 port map( A1 => REGISTERS_0_2_port, A2 => n349, B1 => 
                           REGISTERS_2_2_port, B2 => n312, ZN => n977);
   U1002 : NAND4_X1 port map( A1 => n980, A2 => n979, A3 => n978, A4 => n977, 
                           ZN => n986);
   U1003 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n127_port, B1 =>
                           REGISTERS_15_2_port, B2 => n90, ZN => n984);
   U1004 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n201, B1 => 
                           REGISTERS_11_2_port, B2 => n164, ZN => n983);
   U1005 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n275_port, B1 =>
                           REGISTERS_14_2_port, B2 => n238_port, ZN => n982);
   U1006 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n349, B1 => 
                           REGISTERS_10_2_port, B2 => n312, ZN => n981);
   U1007 : NAND4_X1 port map( A1 => n984, A2 => n983, A3 => n982, A4 => n981, 
                           ZN => n985);
   U1008 : AOI22_X1 port map( A1 => n986, A2 => n27, B1 => n985, B2 => n24, ZN 
                           => n987);
   U1009 : OAI221_X1 port map( B1 => n2271, B2 => n989, C1 => n2269, C2 => n988
                           , A => n987, ZN => N157);
   U1010 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n128_port, B1 =>
                           REGISTERS_23_3_port, B2 => n91, ZN => n993);
   U1011 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n202, B1 => 
                           REGISTERS_19_3_port, B2 => n165, ZN => n992);
   U1012 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n276_port, B1 =>
                           REGISTERS_22_3_port, B2 => n239_port, ZN => n991);
   U1013 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n350, B1 => 
                           REGISTERS_18_3_port, B2 => n313, ZN => n990);
   U1014 : AND4_X1 port map( A1 => n993, A2 => n992, A3 => n991, A4 => n990, ZN
                           => n1010);
   U1015 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n128_port, B1 =>
                           REGISTERS_31_3_port, B2 => n91, ZN => n997);
   U1016 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n202, B1 => 
                           REGISTERS_27_3_port, B2 => n165, ZN => n996);
   U1017 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n276_port, B1 =>
                           REGISTERS_30_3_port, B2 => n239_port, ZN => n995);
   U1018 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n350, B1 => 
                           REGISTERS_26_3_port, B2 => n313, ZN => n994);
   U1019 : AND4_X1 port map( A1 => n997, A2 => n996, A3 => n995, A4 => n994, ZN
                           => n1009);
   U1020 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n128_port, B1 => 
                           REGISTERS_7_3_port, B2 => n91, ZN => n1001);
   U1021 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n202, B1 => 
                           REGISTERS_3_3_port, B2 => n165, ZN => n1000);
   U1022 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n276_port, B1 => 
                           REGISTERS_6_3_port, B2 => n239_port, ZN => n999);
   U1023 : AOI22_X1 port map( A1 => REGISTERS_0_3_port, A2 => n350, B1 => 
                           REGISTERS_2_3_port, B2 => n313, ZN => n998);
   U1024 : NAND4_X1 port map( A1 => n1001, A2 => n1000, A3 => n999, A4 => n998,
                           ZN => n1007);
   U1025 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n128_port, B1 =>
                           REGISTERS_15_3_port, B2 => n91, ZN => n1005);
   U1026 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n202, B1 => 
                           REGISTERS_11_3_port, B2 => n165, ZN => n1004);
   U1027 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n276_port, B1 =>
                           REGISTERS_14_3_port, B2 => n239_port, ZN => n1003);
   U1028 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n350, B1 => 
                           REGISTERS_10_3_port, B2 => n313, ZN => n1002);
   U1029 : NAND4_X1 port map( A1 => n1005, A2 => n1004, A3 => n1003, A4 => 
                           n1002, ZN => n1006);
   U1030 : AOI22_X1 port map( A1 => n1007, A2 => n27, B1 => n1006, B2 => n24, 
                           ZN => n1008);
   U1031 : OAI221_X1 port map( B1 => n2271, B2 => n1010, C1 => n2269, C2 => 
                           n1009, A => n1008, ZN => N156);
   U1032 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n128_port, B1 =>
                           REGISTERS_23_4_port, B2 => n91, ZN => n1014);
   U1033 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n202, B1 => 
                           REGISTERS_19_4_port, B2 => n165, ZN => n1013);
   U1034 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n276_port, B1 =>
                           REGISTERS_22_4_port, B2 => n239_port, ZN => n1012);
   U1035 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n350, B1 => 
                           REGISTERS_18_4_port, B2 => n313, ZN => n1011);
   U1036 : AND4_X1 port map( A1 => n1014, A2 => n1013, A3 => n1012, A4 => n1011
                           , ZN => n1031);
   U1037 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n128_port, B1 =>
                           REGISTERS_31_4_port, B2 => n91, ZN => n1018);
   U1038 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n202, B1 => 
                           REGISTERS_27_4_port, B2 => n165, ZN => n1017);
   U1039 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n276_port, B1 =>
                           REGISTERS_30_4_port, B2 => n239_port, ZN => n1016);
   U1040 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n350, B1 => 
                           REGISTERS_26_4_port, B2 => n313, ZN => n1015);
   U1041 : AND4_X1 port map( A1 => n1018, A2 => n1017, A3 => n1016, A4 => n1015
                           , ZN => n1030);
   U1042 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n128_port, B1 => 
                           REGISTERS_7_4_port, B2 => n91, ZN => n1022);
   U1043 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n202, B1 => 
                           REGISTERS_3_4_port, B2 => n165, ZN => n1021);
   U1044 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n276_port, B1 => 
                           REGISTERS_6_4_port, B2 => n239_port, ZN => n1020);
   U1045 : AOI22_X1 port map( A1 => REGISTERS_0_4_port, A2 => n350, B1 => 
                           REGISTERS_2_4_port, B2 => n313, ZN => n1019);
   U1046 : NAND4_X1 port map( A1 => n1022, A2 => n1021, A3 => n1020, A4 => 
                           n1019, ZN => n1028);
   U1047 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n128_port, B1 =>
                           REGISTERS_15_4_port, B2 => n91, ZN => n1026);
   U1048 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n202, B1 => 
                           REGISTERS_11_4_port, B2 => n165, ZN => n1025);
   U1049 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n276_port, B1 =>
                           REGISTERS_14_4_port, B2 => n239_port, ZN => n1024);
   U1050 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n350, B1 => 
                           REGISTERS_10_4_port, B2 => n313, ZN => n1023);
   U1051 : NAND4_X1 port map( A1 => n1026, A2 => n1025, A3 => n1024, A4 => 
                           n1023, ZN => n1027);
   U1052 : AOI22_X1 port map( A1 => n1028, A2 => n27, B1 => n1027, B2 => n24, 
                           ZN => n1029);
   U1053 : OAI221_X1 port map( B1 => n2271, B2 => n1031, C1 => n2269, C2 => 
                           n1030, A => n1029, ZN => N155);
   U1054 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n128_port, B1 =>
                           REGISTERS_23_5_port, B2 => n91, ZN => n1035);
   U1055 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n202, B1 => 
                           REGISTERS_19_5_port, B2 => n165, ZN => n1034);
   U1056 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n276_port, B1 =>
                           REGISTERS_22_5_port, B2 => n239_port, ZN => n1033);
   U1057 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n350, B1 => 
                           REGISTERS_18_5_port, B2 => n313, ZN => n1032);
   U1058 : AND4_X1 port map( A1 => n1035, A2 => n1034, A3 => n1033, A4 => n1032
                           , ZN => n1052);
   U1059 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n128_port, B1 =>
                           REGISTERS_31_5_port, B2 => n91, ZN => n1039);
   U1060 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n202, B1 => 
                           REGISTERS_27_5_port, B2 => n165, ZN => n1038);
   U1061 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n276_port, B1 =>
                           REGISTERS_30_5_port, B2 => n239_port, ZN => n1037);
   U1062 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n350, B1 => 
                           REGISTERS_26_5_port, B2 => n313, ZN => n1036);
   U1063 : AND4_X1 port map( A1 => n1039, A2 => n1038, A3 => n1037, A4 => n1036
                           , ZN => n1051);
   U1064 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n128_port, B1 => 
                           REGISTERS_7_5_port, B2 => n91, ZN => n1043);
   U1065 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n202, B1 => 
                           REGISTERS_3_5_port, B2 => n165, ZN => n1042);
   U1066 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n276_port, B1 => 
                           REGISTERS_6_5_port, B2 => n239_port, ZN => n1041);
   U1067 : AOI22_X1 port map( A1 => REGISTERS_0_5_port, A2 => n350, B1 => 
                           REGISTERS_2_5_port, B2 => n313, ZN => n1040);
   U1068 : NAND4_X1 port map( A1 => n1043, A2 => n1042, A3 => n1041, A4 => 
                           n1040, ZN => n1049);
   U1069 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n128_port, B1 =>
                           REGISTERS_15_5_port, B2 => n91, ZN => n1047);
   U1070 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n202, B1 => 
                           REGISTERS_11_5_port, B2 => n165, ZN => n1046);
   U1071 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n276_port, B1 =>
                           REGISTERS_14_5_port, B2 => n239_port, ZN => n1045);
   U1072 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n350, B1 => 
                           REGISTERS_10_5_port, B2 => n313, ZN => n1044);
   U1073 : NAND4_X1 port map( A1 => n1047, A2 => n1046, A3 => n1045, A4 => 
                           n1044, ZN => n1048);
   U1074 : AOI22_X1 port map( A1 => n1049, A2 => n27, B1 => n1048, B2 => n24, 
                           ZN => n1050);
   U1075 : OAI221_X1 port map( B1 => n2271, B2 => n1052, C1 => n2269, C2 => 
                           n1051, A => n1050, ZN => N154);
   U1076 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n129_port, B1 =>
                           REGISTERS_23_6_port, B2 => n92, ZN => n1056);
   U1077 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n203, B1 => 
                           REGISTERS_19_6_port, B2 => n166, ZN => n1055);
   U1078 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n277_port, B1 =>
                           REGISTERS_22_6_port, B2 => n240_port, ZN => n1054);
   U1079 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n351, B1 => 
                           REGISTERS_18_6_port, B2 => n314, ZN => n1053);
   U1080 : AND4_X1 port map( A1 => n1056, A2 => n1055, A3 => n1054, A4 => n1053
                           , ZN => n1073);
   U1081 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n129_port, B1 =>
                           REGISTERS_31_6_port, B2 => n92, ZN => n1060);
   U1082 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n203, B1 => 
                           REGISTERS_27_6_port, B2 => n166, ZN => n1059);
   U1083 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n277_port, B1 =>
                           REGISTERS_30_6_port, B2 => n240_port, ZN => n1058);
   U1084 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n351, B1 => 
                           REGISTERS_26_6_port, B2 => n314, ZN => n1057);
   U1085 : AND4_X1 port map( A1 => n1060, A2 => n1059, A3 => n1058, A4 => n1057
                           , ZN => n1072);
   U1086 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n129_port, B1 => 
                           REGISTERS_7_6_port, B2 => n92, ZN => n1064);
   U1087 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n203, B1 => 
                           REGISTERS_3_6_port, B2 => n166, ZN => n1063);
   U1088 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n277_port, B1 => 
                           REGISTERS_6_6_port, B2 => n240_port, ZN => n1062);
   U1089 : AOI22_X1 port map( A1 => REGISTERS_0_6_port, A2 => n351, B1 => 
                           REGISTERS_2_6_port, B2 => n314, ZN => n1061);
   U1090 : NAND4_X1 port map( A1 => n1064, A2 => n1063, A3 => n1062, A4 => 
                           n1061, ZN => n1070);
   U1091 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n129_port, B1 =>
                           REGISTERS_15_6_port, B2 => n92, ZN => n1068);
   U1092 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n203, B1 => 
                           REGISTERS_11_6_port, B2 => n166, ZN => n1067);
   U1093 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n277_port, B1 =>
                           REGISTERS_14_6_port, B2 => n240_port, ZN => n1066);
   U1094 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n351, B1 => 
                           REGISTERS_10_6_port, B2 => n314, ZN => n1065);
   U1095 : NAND4_X1 port map( A1 => n1068, A2 => n1067, A3 => n1066, A4 => 
                           n1065, ZN => n1069);
   U1096 : AOI22_X1 port map( A1 => n1070, A2 => n27, B1 => n1069, B2 => n24, 
                           ZN => n1071);
   U1097 : OAI221_X1 port map( B1 => n2271, B2 => n1073, C1 => n2269, C2 => 
                           n1072, A => n1071, ZN => N153);
   U1098 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n129_port, B1 =>
                           REGISTERS_23_7_port, B2 => n92, ZN => n1077);
   U1099 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n203, B1 => 
                           REGISTERS_19_7_port, B2 => n166, ZN => n1076);
   U1100 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n277_port, B1 =>
                           REGISTERS_22_7_port, B2 => n240_port, ZN => n1075);
   U1101 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n351, B1 => 
                           REGISTERS_18_7_port, B2 => n314, ZN => n1074);
   U1102 : AND4_X1 port map( A1 => n1077, A2 => n1076, A3 => n1075, A4 => n1074
                           , ZN => n1094);
   U1103 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n129_port, B1 =>
                           REGISTERS_31_7_port, B2 => n92, ZN => n1081);
   U1104 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n203, B1 => 
                           REGISTERS_27_7_port, B2 => n166, ZN => n1080);
   U1105 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n277_port, B1 =>
                           REGISTERS_30_7_port, B2 => n240_port, ZN => n1079);
   U1106 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n351, B1 => 
                           REGISTERS_26_7_port, B2 => n314, ZN => n1078);
   U1107 : AND4_X1 port map( A1 => n1081, A2 => n1080, A3 => n1079, A4 => n1078
                           , ZN => n1093);
   U1108 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n129_port, B1 => 
                           REGISTERS_7_7_port, B2 => n92, ZN => n1085);
   U1109 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n203, B1 => 
                           REGISTERS_3_7_port, B2 => n166, ZN => n1084);
   U1110 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n277_port, B1 => 
                           REGISTERS_6_7_port, B2 => n240_port, ZN => n1083);
   U1111 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n351, B1 => 
                           REGISTERS_2_7_port, B2 => n314, ZN => n1082);
   U1112 : NAND4_X1 port map( A1 => n1085, A2 => n1084, A3 => n1083, A4 => 
                           n1082, ZN => n1091);
   U1113 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n129_port, B1 =>
                           REGISTERS_15_7_port, B2 => n92, ZN => n1089);
   U1114 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n203, B1 => 
                           REGISTERS_11_7_port, B2 => n166, ZN => n1088);
   U1115 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n277_port, B1 =>
                           REGISTERS_14_7_port, B2 => n240_port, ZN => n1087);
   U1116 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n351, B1 => 
                           REGISTERS_10_7_port, B2 => n314, ZN => n1086);
   U1117 : NAND4_X1 port map( A1 => n1089, A2 => n1088, A3 => n1087, A4 => 
                           n1086, ZN => n1090);
   U1118 : AOI22_X1 port map( A1 => n1091, A2 => n27, B1 => n1090, B2 => n24, 
                           ZN => n1092);
   U1119 : OAI221_X1 port map( B1 => n2271, B2 => n1094, C1 => n2269, C2 => 
                           n1093, A => n1092, ZN => N152);
   U1120 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n129_port, B1 =>
                           REGISTERS_23_8_port, B2 => n92, ZN => n1098);
   U1121 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n203, B1 => 
                           REGISTERS_19_8_port, B2 => n166, ZN => n1097);
   U1122 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n277_port, B1 =>
                           REGISTERS_22_8_port, B2 => n240_port, ZN => n1096);
   U1123 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n351, B1 => 
                           REGISTERS_18_8_port, B2 => n314, ZN => n1095);
   U1124 : AND4_X1 port map( A1 => n1098, A2 => n1097, A3 => n1096, A4 => n1095
                           , ZN => n1115);
   U1125 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n129_port, B1 =>
                           REGISTERS_31_8_port, B2 => n92, ZN => n1102);
   U1126 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n203, B1 => 
                           REGISTERS_27_8_port, B2 => n166, ZN => n1101);
   U1127 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n277_port, B1 =>
                           REGISTERS_30_8_port, B2 => n240_port, ZN => n1100);
   U1128 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n351, B1 => 
                           REGISTERS_26_8_port, B2 => n314, ZN => n1099);
   U1129 : AND4_X1 port map( A1 => n1102, A2 => n1101, A3 => n1100, A4 => n1099
                           , ZN => n1114);
   U1130 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n129_port, B1 => 
                           REGISTERS_7_8_port, B2 => n92, ZN => n1106);
   U1131 : AOI22_X1 port map( A1 => REGISTERS_1_8_port, A2 => n203, B1 => 
                           REGISTERS_3_8_port, B2 => n166, ZN => n1105);
   U1132 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n277_port, B1 => 
                           REGISTERS_6_8_port, B2 => n240_port, ZN => n1104);
   U1133 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n351, B1 => 
                           REGISTERS_2_8_port, B2 => n314, ZN => n1103);
   U1134 : NAND4_X1 port map( A1 => n1106, A2 => n1105, A3 => n1104, A4 => 
                           n1103, ZN => n1112);
   U1135 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n129_port, B1 =>
                           REGISTERS_15_8_port, B2 => n92, ZN => n1110);
   U1136 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n203, B1 => 
                           REGISTERS_11_8_port, B2 => n166, ZN => n1109);
   U1137 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n277_port, B1 =>
                           REGISTERS_14_8_port, B2 => n240_port, ZN => n1108);
   U1138 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n351, B1 => 
                           REGISTERS_10_8_port, B2 => n314, ZN => n1107);
   U1139 : NAND4_X1 port map( A1 => n1110, A2 => n1109, A3 => n1108, A4 => 
                           n1107, ZN => n1111);
   U1140 : AOI22_X1 port map( A1 => n1112, A2 => n27, B1 => n1111, B2 => n24, 
                           ZN => n1113);
   U1141 : OAI221_X1 port map( B1 => n2271, B2 => n1115, C1 => n2269, C2 => 
                           n1114, A => n1113, ZN => N151);
   U1142 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n130_port, B1 =>
                           REGISTERS_23_9_port, B2 => n93, ZN => n1119);
   U1143 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n204, B1 => 
                           REGISTERS_19_9_port, B2 => n167, ZN => n1118);
   U1144 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n278_port, B1 =>
                           REGISTERS_22_9_port, B2 => n241_port, ZN => n1117);
   U1145 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n352, B1 => 
                           REGISTERS_18_9_port, B2 => n315, ZN => n1116);
   U1146 : AND4_X1 port map( A1 => n1119, A2 => n1118, A3 => n1117, A4 => n1116
                           , ZN => n1136);
   U1147 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n130_port, B1 =>
                           REGISTERS_31_9_port, B2 => n93, ZN => n1123);
   U1148 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n204, B1 => 
                           REGISTERS_27_9_port, B2 => n167, ZN => n1122);
   U1149 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n278_port, B1 =>
                           REGISTERS_30_9_port, B2 => n241_port, ZN => n1121);
   U1150 : AOI22_X1 port map( A1 => REGISTERS_24_9_port, A2 => n352, B1 => 
                           REGISTERS_26_9_port, B2 => n315, ZN => n1120);
   U1151 : AND4_X1 port map( A1 => n1123, A2 => n1122, A3 => n1121, A4 => n1120
                           , ZN => n1135);
   U1152 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n130_port, B1 => 
                           REGISTERS_7_9_port, B2 => n93, ZN => n1127);
   U1153 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n204, B1 => 
                           REGISTERS_3_9_port, B2 => n167, ZN => n1126);
   U1154 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n278_port, B1 => 
                           REGISTERS_6_9_port, B2 => n241_port, ZN => n1125);
   U1155 : AOI22_X1 port map( A1 => REGISTERS_0_9_port, A2 => n352, B1 => 
                           REGISTERS_2_9_port, B2 => n315, ZN => n1124);
   U1156 : NAND4_X1 port map( A1 => n1127, A2 => n1126, A3 => n1125, A4 => 
                           n1124, ZN => n1133);
   U1157 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n130_port, B1 =>
                           REGISTERS_15_9_port, B2 => n93, ZN => n1131);
   U1158 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n204, B1 => 
                           REGISTERS_11_9_port, B2 => n167, ZN => n1130);
   U1159 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n278_port, B1 =>
                           REGISTERS_14_9_port, B2 => n241_port, ZN => n1129);
   U1160 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n352, B1 => 
                           REGISTERS_10_9_port, B2 => n315, ZN => n1128);
   U1161 : NAND4_X1 port map( A1 => n1131, A2 => n1130, A3 => n1129, A4 => 
                           n1128, ZN => n1132);
   U1162 : AOI22_X1 port map( A1 => n1133, A2 => n27, B1 => n1132, B2 => n24, 
                           ZN => n1134);
   U1163 : OAI221_X1 port map( B1 => n2271, B2 => n1136, C1 => n2269, C2 => 
                           n1135, A => n1134, ZN => N150);
   U1164 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n130_port, B1 
                           => REGISTERS_23_10_port, B2 => n93, ZN => n1140);
   U1165 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n204, B1 => 
                           REGISTERS_19_10_port, B2 => n167, ZN => n1139);
   U1166 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n278_port, B1 
                           => REGISTERS_22_10_port, B2 => n241_port, ZN => 
                           n1138);
   U1167 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n352, B1 => 
                           REGISTERS_18_10_port, B2 => n315, ZN => n1137);
   U1168 : AND4_X1 port map( A1 => n1140, A2 => n1139, A3 => n1138, A4 => n1137
                           , ZN => n1157);
   U1169 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n130_port, B1 
                           => REGISTERS_31_10_port, B2 => n93, ZN => n1144);
   U1170 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n204, B1 => 
                           REGISTERS_27_10_port, B2 => n167, ZN => n1143);
   U1171 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n278_port, B1 
                           => REGISTERS_30_10_port, B2 => n241_port, ZN => 
                           n1142);
   U1172 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n352, B1 => 
                           REGISTERS_26_10_port, B2 => n315, ZN => n1141);
   U1173 : AND4_X1 port map( A1 => n1144, A2 => n1143, A3 => n1142, A4 => n1141
                           , ZN => n1156);
   U1174 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n130_port, B1 =>
                           REGISTERS_7_10_port, B2 => n93, ZN => n1148);
   U1175 : AOI22_X1 port map( A1 => REGISTERS_1_10_port, A2 => n204, B1 => 
                           REGISTERS_3_10_port, B2 => n167, ZN => n1147);
   U1176 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n278_port, B1 =>
                           REGISTERS_6_10_port, B2 => n241_port, ZN => n1146);
   U1177 : AOI22_X1 port map( A1 => REGISTERS_0_10_port, A2 => n352, B1 => 
                           REGISTERS_2_10_port, B2 => n315, ZN => n1145);
   U1178 : NAND4_X1 port map( A1 => n1148, A2 => n1147, A3 => n1146, A4 => 
                           n1145, ZN => n1154);
   U1179 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n130_port, B1 
                           => REGISTERS_15_10_port, B2 => n93, ZN => n1152);
   U1180 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n204, B1 => 
                           REGISTERS_11_10_port, B2 => n167, ZN => n1151);
   U1181 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n278_port, B1 
                           => REGISTERS_14_10_port, B2 => n241_port, ZN => 
                           n1150);
   U1182 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n352, B1 => 
                           REGISTERS_10_10_port, B2 => n315, ZN => n1149);
   U1183 : NAND4_X1 port map( A1 => n1152, A2 => n1151, A3 => n1150, A4 => 
                           n1149, ZN => n1153);
   U1184 : AOI22_X1 port map( A1 => n1154, A2 => n27, B1 => n1153, B2 => n24, 
                           ZN => n1155);
   U1185 : OAI221_X1 port map( B1 => n2271, B2 => n1157, C1 => n2269, C2 => 
                           n1156, A => n1155, ZN => N149);
   U1186 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n130_port, B1 
                           => REGISTERS_23_11_port, B2 => n93, ZN => n1161);
   U1187 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n204, B1 => 
                           REGISTERS_19_11_port, B2 => n167, ZN => n1160);
   U1188 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n278_port, B1 
                           => REGISTERS_22_11_port, B2 => n241_port, ZN => 
                           n1159);
   U1189 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n352, B1 => 
                           REGISTERS_18_11_port, B2 => n315, ZN => n1158);
   U1190 : AND4_X1 port map( A1 => n1161, A2 => n1160, A3 => n1159, A4 => n1158
                           , ZN => n1178);
   U1191 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n130_port, B1 
                           => REGISTERS_31_11_port, B2 => n93, ZN => n1165);
   U1192 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n204, B1 => 
                           REGISTERS_27_11_port, B2 => n167, ZN => n1164);
   U1193 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n278_port, B1 
                           => REGISTERS_30_11_port, B2 => n241_port, ZN => 
                           n1163);
   U1194 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n352, B1 => 
                           REGISTERS_26_11_port, B2 => n315, ZN => n1162);
   U1195 : AND4_X1 port map( A1 => n1165, A2 => n1164, A3 => n1163, A4 => n1162
                           , ZN => n1177);
   U1196 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n130_port, B1 =>
                           REGISTERS_7_11_port, B2 => n93, ZN => n1169);
   U1197 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n204, B1 => 
                           REGISTERS_3_11_port, B2 => n167, ZN => n1168);
   U1198 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n278_port, B1 =>
                           REGISTERS_6_11_port, B2 => n241_port, ZN => n1167);
   U1199 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n352, B1 => 
                           REGISTERS_2_11_port, B2 => n315, ZN => n1166);
   U1200 : NAND4_X1 port map( A1 => n1169, A2 => n1168, A3 => n1167, A4 => 
                           n1166, ZN => n1175);
   U1201 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n130_port, B1 
                           => REGISTERS_15_11_port, B2 => n93, ZN => n1173);
   U1202 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n204, B1 => 
                           REGISTERS_11_11_port, B2 => n167, ZN => n1172);
   U1203 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n278_port, B1 
                           => REGISTERS_14_11_port, B2 => n241_port, ZN => 
                           n1171);
   U1204 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n352, B1 => 
                           REGISTERS_10_11_port, B2 => n315, ZN => n1170);
   U1205 : NAND4_X1 port map( A1 => n1173, A2 => n1172, A3 => n1171, A4 => 
                           n1170, ZN => n1174);
   U1206 : AOI22_X1 port map( A1 => n1175, A2 => n27, B1 => n1174, B2 => n24, 
                           ZN => n1176);
   U1207 : OAI221_X1 port map( B1 => n2271, B2 => n1178, C1 => n2269, C2 => 
                           n1177, A => n1176, ZN => N148);
   U1208 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n131_port, B1 
                           => REGISTERS_23_12_port, B2 => n94, ZN => n1182);
   U1209 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n205, B1 => 
                           REGISTERS_19_12_port, B2 => n168, ZN => n1181);
   U1210 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n279_port, B1 
                           => REGISTERS_22_12_port, B2 => n242_port, ZN => 
                           n1180);
   U1211 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n353, B1 => 
                           REGISTERS_18_12_port, B2 => n316, ZN => n1179);
   U1212 : AND4_X1 port map( A1 => n1182, A2 => n1181, A3 => n1180, A4 => n1179
                           , ZN => n1199);
   U1213 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n131_port, B1 
                           => REGISTERS_31_12_port, B2 => n94, ZN => n1186);
   U1214 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n205, B1 => 
                           REGISTERS_27_12_port, B2 => n168, ZN => n1185);
   U1215 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n279_port, B1 
                           => REGISTERS_30_12_port, B2 => n242_port, ZN => 
                           n1184);
   U1216 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n353, B1 => 
                           REGISTERS_26_12_port, B2 => n316, ZN => n1183);
   U1217 : AND4_X1 port map( A1 => n1186, A2 => n1185, A3 => n1184, A4 => n1183
                           , ZN => n1198);
   U1218 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n131_port, B1 =>
                           REGISTERS_7_12_port, B2 => n94, ZN => n1190);
   U1219 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n205, B1 => 
                           REGISTERS_3_12_port, B2 => n168, ZN => n1189);
   U1220 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n279_port, B1 =>
                           REGISTERS_6_12_port, B2 => n242_port, ZN => n1188);
   U1221 : AOI22_X1 port map( A1 => REGISTERS_0_12_port, A2 => n353, B1 => 
                           REGISTERS_2_12_port, B2 => n316, ZN => n1187);
   U1222 : NAND4_X1 port map( A1 => n1190, A2 => n1189, A3 => n1188, A4 => 
                           n1187, ZN => n1196);
   U1223 : AOI22_X1 port map( A1 => REGISTERS_13_12_port, A2 => n131_port, B1 
                           => REGISTERS_15_12_port, B2 => n94, ZN => n1194);
   U1224 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n205, B1 => 
                           REGISTERS_11_12_port, B2 => n168, ZN => n1193);
   U1225 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n279_port, B1 
                           => REGISTERS_14_12_port, B2 => n242_port, ZN => 
                           n1192);
   U1226 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n353, B1 => 
                           REGISTERS_10_12_port, B2 => n316, ZN => n1191);
   U1227 : NAND4_X1 port map( A1 => n1194, A2 => n1193, A3 => n1192, A4 => 
                           n1191, ZN => n1195);
   U1228 : AOI22_X1 port map( A1 => n1196, A2 => n27, B1 => n1195, B2 => n24, 
                           ZN => n1197);
   U1229 : OAI221_X1 port map( B1 => n2271, B2 => n1199, C1 => n2269, C2 => 
                           n1198, A => n1197, ZN => N147);
   U1230 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n131_port, B1 
                           => REGISTERS_23_13_port, B2 => n94, ZN => n1203);
   U1231 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n205, B1 => 
                           REGISTERS_19_13_port, B2 => n168, ZN => n1202);
   U1232 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n279_port, B1 
                           => REGISTERS_22_13_port, B2 => n242_port, ZN => 
                           n1201);
   U1233 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n353, B1 => 
                           REGISTERS_18_13_port, B2 => n316, ZN => n1200);
   U1234 : AND4_X1 port map( A1 => n1203, A2 => n1202, A3 => n1201, A4 => n1200
                           , ZN => n1220);
   U1235 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n131_port, B1 
                           => REGISTERS_31_13_port, B2 => n94, ZN => n1207);
   U1236 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n205, B1 => 
                           REGISTERS_27_13_port, B2 => n168, ZN => n1206);
   U1237 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n279_port, B1 
                           => REGISTERS_30_13_port, B2 => n242_port, ZN => 
                           n1205);
   U1238 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n353, B1 => 
                           REGISTERS_26_13_port, B2 => n316, ZN => n1204);
   U1239 : AND4_X1 port map( A1 => n1207, A2 => n1206, A3 => n1205, A4 => n1204
                           , ZN => n1219);
   U1240 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n131_port, B1 =>
                           REGISTERS_7_13_port, B2 => n94, ZN => n1211);
   U1241 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n205, B1 => 
                           REGISTERS_3_13_port, B2 => n168, ZN => n1210);
   U1242 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n279_port, B1 =>
                           REGISTERS_6_13_port, B2 => n242_port, ZN => n1209);
   U1243 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n353, B1 => 
                           REGISTERS_2_13_port, B2 => n316, ZN => n1208);
   U1244 : NAND4_X1 port map( A1 => n1211, A2 => n1210, A3 => n1209, A4 => 
                           n1208, ZN => n1217);
   U1245 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n131_port, B1 
                           => REGISTERS_15_13_port, B2 => n94, ZN => n1215);
   U1246 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n205, B1 => 
                           REGISTERS_11_13_port, B2 => n168, ZN => n1214);
   U1247 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n279_port, B1 
                           => REGISTERS_14_13_port, B2 => n242_port, ZN => 
                           n1213);
   U1248 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n353, B1 => 
                           REGISTERS_10_13_port, B2 => n316, ZN => n1212);
   U1249 : NAND4_X1 port map( A1 => n1215, A2 => n1214, A3 => n1213, A4 => 
                           n1212, ZN => n1216);
   U1250 : AOI22_X1 port map( A1 => n1217, A2 => n27, B1 => n1216, B2 => n24, 
                           ZN => n1218);
   U1251 : OAI221_X1 port map( B1 => n2271, B2 => n1220, C1 => n2269, C2 => 
                           n1219, A => n1218, ZN => N146);
   U1252 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n131_port, B1 
                           => REGISTERS_23_14_port, B2 => n94, ZN => n1224);
   U1253 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n205, B1 => 
                           REGISTERS_19_14_port, B2 => n168, ZN => n1223);
   U1254 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n279_port, B1 
                           => REGISTERS_22_14_port, B2 => n242_port, ZN => 
                           n1222);
   U1255 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n353, B1 => 
                           REGISTERS_18_14_port, B2 => n316, ZN => n1221);
   U1256 : AND4_X1 port map( A1 => n1224, A2 => n1223, A3 => n1222, A4 => n1221
                           , ZN => n1241);
   U1257 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n131_port, B1 
                           => REGISTERS_31_14_port, B2 => n94, ZN => n1228);
   U1258 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n205, B1 => 
                           REGISTERS_27_14_port, B2 => n168, ZN => n1227);
   U1259 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n279_port, B1 
                           => REGISTERS_30_14_port, B2 => n242_port, ZN => 
                           n1226);
   U1260 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n353, B1 => 
                           REGISTERS_26_14_port, B2 => n316, ZN => n1225);
   U1261 : AND4_X1 port map( A1 => n1228, A2 => n1227, A3 => n1226, A4 => n1225
                           , ZN => n1240);
   U1262 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n131_port, B1 =>
                           REGISTERS_7_14_port, B2 => n94, ZN => n1232);
   U1263 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n205, B1 => 
                           REGISTERS_3_14_port, B2 => n168, ZN => n1231);
   U1264 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n279_port, B1 =>
                           REGISTERS_6_14_port, B2 => n242_port, ZN => n1230);
   U1265 : AOI22_X1 port map( A1 => REGISTERS_0_14_port, A2 => n353, B1 => 
                           REGISTERS_2_14_port, B2 => n316, ZN => n1229);
   U1266 : NAND4_X1 port map( A1 => n1232, A2 => n1231, A3 => n1230, A4 => 
                           n1229, ZN => n1238);
   U1267 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n131_port, B1 
                           => REGISTERS_15_14_port, B2 => n94, ZN => n1236);
   U1268 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n205, B1 => 
                           REGISTERS_11_14_port, B2 => n168, ZN => n1235);
   U1269 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n279_port, B1 
                           => REGISTERS_14_14_port, B2 => n242_port, ZN => 
                           n1234);
   U1270 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n353, B1 => 
                           REGISTERS_10_14_port, B2 => n316, ZN => n1233);
   U1271 : NAND4_X1 port map( A1 => n1236, A2 => n1235, A3 => n1234, A4 => 
                           n1233, ZN => n1237);
   U1272 : AOI22_X1 port map( A1 => n1238, A2 => n27, B1 => n1237, B2 => n24, 
                           ZN => n1239);
   U1273 : OAI221_X1 port map( B1 => n2271, B2 => n1241, C1 => n2269, C2 => 
                           n1240, A => n1239, ZN => N145);
   U1274 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n132_port, B1 
                           => REGISTERS_23_15_port, B2 => n95, ZN => n1245);
   U1275 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n206, B1 => 
                           REGISTERS_19_15_port, B2 => n169, ZN => n1244);
   U1276 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n280_port, B1 
                           => REGISTERS_22_15_port, B2 => n243_port, ZN => 
                           n1243);
   U1277 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n354, B1 => 
                           REGISTERS_18_15_port, B2 => n317, ZN => n1242);
   U1278 : AND4_X1 port map( A1 => n1245, A2 => n1244, A3 => n1243, A4 => n1242
                           , ZN => n1262);
   U1279 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n132_port, B1 
                           => REGISTERS_31_15_port, B2 => n95, ZN => n1249);
   U1280 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n206, B1 => 
                           REGISTERS_27_15_port, B2 => n169, ZN => n1248);
   U1281 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n280_port, B1 
                           => REGISTERS_30_15_port, B2 => n243_port, ZN => 
                           n1247);
   U1282 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n354, B1 => 
                           REGISTERS_26_15_port, B2 => n317, ZN => n1246);
   U1283 : AND4_X1 port map( A1 => n1249, A2 => n1248, A3 => n1247, A4 => n1246
                           , ZN => n1261);
   U1284 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n132_port, B1 =>
                           REGISTERS_7_15_port, B2 => n95, ZN => n1253);
   U1285 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n206, B1 => 
                           REGISTERS_3_15_port, B2 => n169, ZN => n1252);
   U1286 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n280_port, B1 =>
                           REGISTERS_6_15_port, B2 => n243_port, ZN => n1251);
   U1287 : AOI22_X1 port map( A1 => REGISTERS_0_15_port, A2 => n354, B1 => 
                           REGISTERS_2_15_port, B2 => n317, ZN => n1250);
   U1288 : NAND4_X1 port map( A1 => n1253, A2 => n1252, A3 => n1251, A4 => 
                           n1250, ZN => n1259);
   U1289 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n132_port, B1 
                           => REGISTERS_15_15_port, B2 => n95, ZN => n1257);
   U1290 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n206, B1 => 
                           REGISTERS_11_15_port, B2 => n169, ZN => n1256);
   U1291 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n280_port, B1 
                           => REGISTERS_14_15_port, B2 => n243_port, ZN => 
                           n1255);
   U1292 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n354, B1 => 
                           REGISTERS_10_15_port, B2 => n317, ZN => n1254);
   U1293 : NAND4_X1 port map( A1 => n1257, A2 => n1256, A3 => n1255, A4 => 
                           n1254, ZN => n1258);
   U1294 : AOI22_X1 port map( A1 => n1259, A2 => n27, B1 => n1258, B2 => n24, 
                           ZN => n1260);
   U1295 : OAI221_X1 port map( B1 => n2271, B2 => n1262, C1 => n2269, C2 => 
                           n1261, A => n1260, ZN => N144);
   U1296 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n132_port, B1 
                           => REGISTERS_23_16_port, B2 => n95, ZN => n1266);
   U1297 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n206, B1 => 
                           REGISTERS_19_16_port, B2 => n169, ZN => n1265);
   U1298 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n280_port, B1 
                           => REGISTERS_22_16_port, B2 => n243_port, ZN => 
                           n1264);
   U1299 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n354, B1 => 
                           REGISTERS_18_16_port, B2 => n317, ZN => n1263);
   U1300 : AND4_X1 port map( A1 => n1266, A2 => n1265, A3 => n1264, A4 => n1263
                           , ZN => n1283);
   U1301 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n132_port, B1 
                           => REGISTERS_31_16_port, B2 => n95, ZN => n1270);
   U1302 : AOI22_X1 port map( A1 => REGISTERS_25_16_port, A2 => n206, B1 => 
                           REGISTERS_27_16_port, B2 => n169, ZN => n1269);
   U1303 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n280_port, B1 
                           => REGISTERS_30_16_port, B2 => n243_port, ZN => 
                           n1268);
   U1304 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n354, B1 => 
                           REGISTERS_26_16_port, B2 => n317, ZN => n1267);
   U1305 : AND4_X1 port map( A1 => n1270, A2 => n1269, A3 => n1268, A4 => n1267
                           , ZN => n1282);
   U1306 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n132_port, B1 =>
                           REGISTERS_7_16_port, B2 => n95, ZN => n1274);
   U1307 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n206, B1 => 
                           REGISTERS_3_16_port, B2 => n169, ZN => n1273);
   U1308 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n280_port, B1 =>
                           REGISTERS_6_16_port, B2 => n243_port, ZN => n1272);
   U1309 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n354, B1 => 
                           REGISTERS_2_16_port, B2 => n317, ZN => n1271);
   U1310 : NAND4_X1 port map( A1 => n1274, A2 => n1273, A3 => n1272, A4 => 
                           n1271, ZN => n1280);
   U1311 : AOI22_X1 port map( A1 => REGISTERS_13_16_port, A2 => n132_port, B1 
                           => REGISTERS_15_16_port, B2 => n95, ZN => n1278);
   U1312 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n206, B1 => 
                           REGISTERS_11_16_port, B2 => n169, ZN => n1277);
   U1313 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n280_port, B1 
                           => REGISTERS_14_16_port, B2 => n243_port, ZN => 
                           n1276);
   U1314 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n354, B1 => 
                           REGISTERS_10_16_port, B2 => n317, ZN => n1275);
   U1315 : NAND4_X1 port map( A1 => n1278, A2 => n1277, A3 => n1276, A4 => 
                           n1275, ZN => n1279);
   U1316 : AOI22_X1 port map( A1 => n1280, A2 => n27, B1 => n1279, B2 => n24, 
                           ZN => n1281);
   U1317 : OAI221_X1 port map( B1 => n2271, B2 => n1283, C1 => n2269, C2 => 
                           n1282, A => n1281, ZN => N143);
   U1318 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n132_port, B1 
                           => REGISTERS_23_17_port, B2 => n95, ZN => n1287);
   U1319 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n206, B1 => 
                           REGISTERS_19_17_port, B2 => n169, ZN => n1286);
   U1320 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n280_port, B1 
                           => REGISTERS_22_17_port, B2 => n243_port, ZN => 
                           n1285);
   U1321 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n354, B1 => 
                           REGISTERS_18_17_port, B2 => n317, ZN => n1284);
   U1322 : AND4_X1 port map( A1 => n1287, A2 => n1286, A3 => n1285, A4 => n1284
                           , ZN => n1304);
   U1323 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n132_port, B1 
                           => REGISTERS_31_17_port, B2 => n95, ZN => n1291);
   U1324 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n206, B1 => 
                           REGISTERS_27_17_port, B2 => n169, ZN => n1290);
   U1325 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n280_port, B1 
                           => REGISTERS_30_17_port, B2 => n243_port, ZN => 
                           n1289);
   U1326 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n354, B1 => 
                           REGISTERS_26_17_port, B2 => n317, ZN => n1288);
   U1327 : AND4_X1 port map( A1 => n1291, A2 => n1290, A3 => n1289, A4 => n1288
                           , ZN => n1303);
   U1328 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n132_port, B1 =>
                           REGISTERS_7_17_port, B2 => n95, ZN => n1295);
   U1329 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n206, B1 => 
                           REGISTERS_3_17_port, B2 => n169, ZN => n1294);
   U1330 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n280_port, B1 =>
                           REGISTERS_6_17_port, B2 => n243_port, ZN => n1293);
   U1331 : AOI22_X1 port map( A1 => REGISTERS_0_17_port, A2 => n354, B1 => 
                           REGISTERS_2_17_port, B2 => n317, ZN => n1292);
   U1332 : NAND4_X1 port map( A1 => n1295, A2 => n1294, A3 => n1293, A4 => 
                           n1292, ZN => n1301);
   U1333 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n132_port, B1 
                           => REGISTERS_15_17_port, B2 => n95, ZN => n1299);
   U1334 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n206, B1 => 
                           REGISTERS_11_17_port, B2 => n169, ZN => n1298);
   U1335 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n280_port, B1 
                           => REGISTERS_14_17_port, B2 => n243_port, ZN => 
                           n1297);
   U1336 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n354, B1 => 
                           REGISTERS_10_17_port, B2 => n317, ZN => n1296);
   U1337 : NAND4_X1 port map( A1 => n1299, A2 => n1298, A3 => n1297, A4 => 
                           n1296, ZN => n1300);
   U1338 : AOI22_X1 port map( A1 => n1301, A2 => n27, B1 => n1300, B2 => n24, 
                           ZN => n1302);
   U1339 : OAI221_X1 port map( B1 => n2271, B2 => n1304, C1 => n2269, C2 => 
                           n1303, A => n1302, ZN => N142);
   U1340 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n133_port, B1 
                           => REGISTERS_23_18_port, B2 => n96_port, ZN => n1308
                           );
   U1341 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n207, B1 => 
                           REGISTERS_19_18_port, B2 => n170, ZN => n1307);
   U1342 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n281_port, B1 
                           => REGISTERS_22_18_port, B2 => n244_port, ZN => 
                           n1306);
   U1343 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n355, B1 => 
                           REGISTERS_18_18_port, B2 => n318, ZN => n1305);
   U1344 : AND4_X1 port map( A1 => n1308, A2 => n1307, A3 => n1306, A4 => n1305
                           , ZN => n1325);
   U1345 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n133_port, B1 
                           => REGISTERS_31_18_port, B2 => n96_port, ZN => n1312
                           );
   U1346 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n207, B1 => 
                           REGISTERS_27_18_port, B2 => n170, ZN => n1311);
   U1347 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n281_port, B1 
                           => REGISTERS_30_18_port, B2 => n244_port, ZN => 
                           n1310);
   U1348 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n355, B1 => 
                           REGISTERS_26_18_port, B2 => n318, ZN => n1309);
   U1349 : AND4_X1 port map( A1 => n1312, A2 => n1311, A3 => n1310, A4 => n1309
                           , ZN => n1324);
   U1350 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n133_port, B1 =>
                           REGISTERS_7_18_port, B2 => n96_port, ZN => n1316);
   U1351 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n207, B1 => 
                           REGISTERS_3_18_port, B2 => n170, ZN => n1315);
   U1352 : AOI22_X1 port map( A1 => REGISTERS_4_18_port, A2 => n281_port, B1 =>
                           REGISTERS_6_18_port, B2 => n244_port, ZN => n1314);
   U1353 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n355, B1 => 
                           REGISTERS_2_18_port, B2 => n318, ZN => n1313);
   U1354 : NAND4_X1 port map( A1 => n1316, A2 => n1315, A3 => n1314, A4 => 
                           n1313, ZN => n1322);
   U1355 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n133_port, B1 
                           => REGISTERS_15_18_port, B2 => n96_port, ZN => n1320
                           );
   U1356 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n207, B1 => 
                           REGISTERS_11_18_port, B2 => n170, ZN => n1319);
   U1357 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n281_port, B1 
                           => REGISTERS_14_18_port, B2 => n244_port, ZN => 
                           n1318);
   U1358 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n355, B1 => 
                           REGISTERS_10_18_port, B2 => n318, ZN => n1317);
   U1359 : NAND4_X1 port map( A1 => n1320, A2 => n1319, A3 => n1318, A4 => 
                           n1317, ZN => n1321);
   U1360 : AOI22_X1 port map( A1 => n1322, A2 => n27, B1 => n1321, B2 => n24, 
                           ZN => n1323);
   U1361 : OAI221_X1 port map( B1 => n2271, B2 => n1325, C1 => n2269, C2 => 
                           n1324, A => n1323, ZN => N141);
   U1362 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n133_port, B1 
                           => REGISTERS_23_19_port, B2 => n96_port, ZN => n1329
                           );
   U1363 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n207, B1 => 
                           REGISTERS_19_19_port, B2 => n170, ZN => n1328);
   U1364 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n281_port, B1 
                           => REGISTERS_22_19_port, B2 => n244_port, ZN => 
                           n1327);
   U1365 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n355, B1 => 
                           REGISTERS_18_19_port, B2 => n318, ZN => n1326);
   U1366 : AND4_X1 port map( A1 => n1329, A2 => n1328, A3 => n1327, A4 => n1326
                           , ZN => n1346);
   U1367 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n133_port, B1 
                           => REGISTERS_31_19_port, B2 => n96_port, ZN => n1333
                           );
   U1368 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n207, B1 => 
                           REGISTERS_27_19_port, B2 => n170, ZN => n1332);
   U1369 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n281_port, B1 
                           => REGISTERS_30_19_port, B2 => n244_port, ZN => 
                           n1331);
   U1370 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n355, B1 => 
                           REGISTERS_26_19_port, B2 => n318, ZN => n1330);
   U1371 : AND4_X1 port map( A1 => n1333, A2 => n1332, A3 => n1331, A4 => n1330
                           , ZN => n1345);
   U1372 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n133_port, B1 =>
                           REGISTERS_7_19_port, B2 => n96_port, ZN => n1337);
   U1373 : AOI22_X1 port map( A1 => REGISTERS_1_19_port, A2 => n207, B1 => 
                           REGISTERS_3_19_port, B2 => n170, ZN => n1336);
   U1374 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n281_port, B1 =>
                           REGISTERS_6_19_port, B2 => n244_port, ZN => n1335);
   U1375 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n355, B1 => 
                           REGISTERS_2_19_port, B2 => n318, ZN => n1334);
   U1376 : NAND4_X1 port map( A1 => n1337, A2 => n1336, A3 => n1335, A4 => 
                           n1334, ZN => n1343);
   U1377 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n133_port, B1 
                           => REGISTERS_15_19_port, B2 => n96_port, ZN => n1341
                           );
   U1378 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n207, B1 => 
                           REGISTERS_11_19_port, B2 => n170, ZN => n1340);
   U1379 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n281_port, B1 
                           => REGISTERS_14_19_port, B2 => n244_port, ZN => 
                           n1339);
   U1380 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n355, B1 => 
                           REGISTERS_10_19_port, B2 => n318, ZN => n1338);
   U1381 : NAND4_X1 port map( A1 => n1341, A2 => n1340, A3 => n1339, A4 => 
                           n1338, ZN => n1342);
   U1382 : AOI22_X1 port map( A1 => n1343, A2 => n27, B1 => n1342, B2 => n24, 
                           ZN => n1344);
   U1383 : OAI221_X1 port map( B1 => n2271, B2 => n1346, C1 => n2269, C2 => 
                           n1345, A => n1344, ZN => N140);
   U1384 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n133_port, B1 
                           => REGISTERS_23_20_port, B2 => n96_port, ZN => n1350
                           );
   U1385 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n207, B1 => 
                           REGISTERS_19_20_port, B2 => n170, ZN => n1349);
   U1386 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n281_port, B1 
                           => REGISTERS_22_20_port, B2 => n244_port, ZN => 
                           n1348);
   U1387 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n355, B1 => 
                           REGISTERS_18_20_port, B2 => n318, ZN => n1347);
   U1388 : AND4_X1 port map( A1 => n1350, A2 => n1349, A3 => n1348, A4 => n1347
                           , ZN => n1367);
   U1389 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n133_port, B1 
                           => REGISTERS_31_20_port, B2 => n96_port, ZN => n1354
                           );
   U1390 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n207, B1 => 
                           REGISTERS_27_20_port, B2 => n170, ZN => n1353);
   U1391 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n281_port, B1 
                           => REGISTERS_30_20_port, B2 => n244_port, ZN => 
                           n1352);
   U1392 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n355, B1 => 
                           REGISTERS_26_20_port, B2 => n318, ZN => n1351);
   U1393 : AND4_X1 port map( A1 => n1354, A2 => n1353, A3 => n1352, A4 => n1351
                           , ZN => n1366);
   U1394 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n133_port, B1 =>
                           REGISTERS_7_20_port, B2 => n96_port, ZN => n1358);
   U1395 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n207, B1 => 
                           REGISTERS_3_20_port, B2 => n170, ZN => n1357);
   U1396 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n281_port, B1 =>
                           REGISTERS_6_20_port, B2 => n244_port, ZN => n1356);
   U1397 : AOI22_X1 port map( A1 => REGISTERS_0_20_port, A2 => n355, B1 => 
                           REGISTERS_2_20_port, B2 => n318, ZN => n1355);
   U1398 : NAND4_X1 port map( A1 => n1358, A2 => n1357, A3 => n1356, A4 => 
                           n1355, ZN => n1364);
   U1399 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n133_port, B1 
                           => REGISTERS_15_20_port, B2 => n96_port, ZN => n1362
                           );
   U1400 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n207, B1 => 
                           REGISTERS_11_20_port, B2 => n170, ZN => n1361);
   U1401 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n281_port, B1 
                           => REGISTERS_14_20_port, B2 => n244_port, ZN => 
                           n1360);
   U1402 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n355, B1 => 
                           REGISTERS_10_20_port, B2 => n318, ZN => n1359);
   U1403 : NAND4_X1 port map( A1 => n1362, A2 => n1361, A3 => n1360, A4 => 
                           n1359, ZN => n1363);
   U1404 : AOI22_X1 port map( A1 => n1364, A2 => n27, B1 => n1363, B2 => n24, 
                           ZN => n1365);
   U1405 : OAI221_X1 port map( B1 => n2271, B2 => n1367, C1 => n2269, C2 => 
                           n1366, A => n1365, ZN => N139);
   U1406 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n134_port, B1 
                           => REGISTERS_23_21_port, B2 => n97_port, ZN => n1371
                           );
   U1407 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n208, B1 => 
                           REGISTERS_19_21_port, B2 => n171, ZN => n1370);
   U1408 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n282_port, B1 
                           => REGISTERS_22_21_port, B2 => n245_port, ZN => 
                           n1369);
   U1409 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n356, B1 => 
                           REGISTERS_18_21_port, B2 => n319, ZN => n1368);
   U1410 : AND4_X1 port map( A1 => n1371, A2 => n1370, A3 => n1369, A4 => n1368
                           , ZN => n1388);
   U1411 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n134_port, B1 
                           => REGISTERS_31_21_port, B2 => n97_port, ZN => n1375
                           );
   U1412 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n208, B1 => 
                           REGISTERS_27_21_port, B2 => n171, ZN => n1374);
   U1413 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n282_port, B1 
                           => REGISTERS_30_21_port, B2 => n245_port, ZN => 
                           n1373);
   U1414 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n356, B1 => 
                           REGISTERS_26_21_port, B2 => n319, ZN => n1372);
   U1415 : AND4_X1 port map( A1 => n1375, A2 => n1374, A3 => n1373, A4 => n1372
                           , ZN => n1387);
   U1416 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n134_port, B1 =>
                           REGISTERS_7_21_port, B2 => n97_port, ZN => n1379);
   U1417 : AOI22_X1 port map( A1 => REGISTERS_1_21_port, A2 => n208, B1 => 
                           REGISTERS_3_21_port, B2 => n171, ZN => n1378);
   U1418 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n282_port, B1 =>
                           REGISTERS_6_21_port, B2 => n245_port, ZN => n1377);
   U1419 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n356, B1 => 
                           REGISTERS_2_21_port, B2 => n319, ZN => n1376);
   U1420 : NAND4_X1 port map( A1 => n1379, A2 => n1378, A3 => n1377, A4 => 
                           n1376, ZN => n1385);
   U1421 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n134_port, B1 
                           => REGISTERS_15_21_port, B2 => n97_port, ZN => n1383
                           );
   U1422 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n208, B1 => 
                           REGISTERS_11_21_port, B2 => n171, ZN => n1382);
   U1423 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n282_port, B1 
                           => REGISTERS_14_21_port, B2 => n245_port, ZN => 
                           n1381);
   U1424 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n356, B1 => 
                           REGISTERS_10_21_port, B2 => n319, ZN => n1380);
   U1425 : NAND4_X1 port map( A1 => n1383, A2 => n1382, A3 => n1381, A4 => 
                           n1380, ZN => n1384);
   U1426 : AOI22_X1 port map( A1 => n1385, A2 => n27, B1 => n1384, B2 => n24, 
                           ZN => n1386);
   U1427 : OAI221_X1 port map( B1 => n2271, B2 => n1388, C1 => n2269, C2 => 
                           n1387, A => n1386, ZN => N138);
   U1428 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n134_port, B1 
                           => REGISTERS_23_22_port, B2 => n97_port, ZN => n1392
                           );
   U1429 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n208, B1 => 
                           REGISTERS_19_22_port, B2 => n171, ZN => n1391);
   U1430 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n282_port, B1 
                           => REGISTERS_22_22_port, B2 => n245_port, ZN => 
                           n1390);
   U1431 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n356, B1 => 
                           REGISTERS_18_22_port, B2 => n319, ZN => n1389);
   U1432 : AND4_X1 port map( A1 => n1392, A2 => n1391, A3 => n1390, A4 => n1389
                           , ZN => n1409);
   U1433 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n134_port, B1 
                           => REGISTERS_31_22_port, B2 => n97_port, ZN => n1396
                           );
   U1434 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n208, B1 => 
                           REGISTERS_27_22_port, B2 => n171, ZN => n1395);
   U1435 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n282_port, B1 
                           => REGISTERS_30_22_port, B2 => n245_port, ZN => 
                           n1394);
   U1436 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n356, B1 => 
                           REGISTERS_26_22_port, B2 => n319, ZN => n1393);
   U1437 : AND4_X1 port map( A1 => n1396, A2 => n1395, A3 => n1394, A4 => n1393
                           , ZN => n1408);
   U1438 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n134_port, B1 =>
                           REGISTERS_7_22_port, B2 => n97_port, ZN => n1400);
   U1439 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n208, B1 => 
                           REGISTERS_3_22_port, B2 => n171, ZN => n1399);
   U1440 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n282_port, B1 =>
                           REGISTERS_6_22_port, B2 => n245_port, ZN => n1398);
   U1441 : AOI22_X1 port map( A1 => REGISTERS_0_22_port, A2 => n356, B1 => 
                           REGISTERS_2_22_port, B2 => n319, ZN => n1397);
   U1442 : NAND4_X1 port map( A1 => n1400, A2 => n1399, A3 => n1398, A4 => 
                           n1397, ZN => n1406);
   U1443 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n134_port, B1 
                           => REGISTERS_15_22_port, B2 => n97_port, ZN => n1404
                           );
   U1444 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n208, B1 => 
                           REGISTERS_11_22_port, B2 => n171, ZN => n1403);
   U1445 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n282_port, B1 
                           => REGISTERS_14_22_port, B2 => n245_port, ZN => 
                           n1402);
   U1446 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n356, B1 => 
                           REGISTERS_10_22_port, B2 => n319, ZN => n1401);
   U1447 : NAND4_X1 port map( A1 => n1404, A2 => n1403, A3 => n1402, A4 => 
                           n1401, ZN => n1405);
   U1448 : AOI22_X1 port map( A1 => n1406, A2 => n27, B1 => n1405, B2 => n24, 
                           ZN => n1407);
   U1449 : OAI221_X1 port map( B1 => n2271, B2 => n1409, C1 => n2269, C2 => 
                           n1408, A => n1407, ZN => N137);
   U1450 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n134_port, B1 
                           => REGISTERS_23_23_port, B2 => n97_port, ZN => n1413
                           );
   U1451 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n208, B1 => 
                           REGISTERS_19_23_port, B2 => n171, ZN => n1412);
   U1452 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n282_port, B1 
                           => REGISTERS_22_23_port, B2 => n245_port, ZN => 
                           n1411);
   U1453 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n356, B1 => 
                           REGISTERS_18_23_port, B2 => n319, ZN => n1410);
   U1454 : AND4_X1 port map( A1 => n1413, A2 => n1412, A3 => n1411, A4 => n1410
                           , ZN => n1430);
   U1455 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n134_port, B1 
                           => REGISTERS_31_23_port, B2 => n97_port, ZN => n1417
                           );
   U1456 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n208, B1 => 
                           REGISTERS_27_23_port, B2 => n171, ZN => n1416);
   U1457 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n282_port, B1 
                           => REGISTERS_30_23_port, B2 => n245_port, ZN => 
                           n1415);
   U1458 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n356, B1 => 
                           REGISTERS_26_23_port, B2 => n319, ZN => n1414);
   U1459 : AND4_X1 port map( A1 => n1417, A2 => n1416, A3 => n1415, A4 => n1414
                           , ZN => n1429);
   U1460 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n134_port, B1 =>
                           REGISTERS_7_23_port, B2 => n97_port, ZN => n1421);
   U1461 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n208, B1 => 
                           REGISTERS_3_23_port, B2 => n171, ZN => n1420);
   U1462 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n282_port, B1 =>
                           REGISTERS_6_23_port, B2 => n245_port, ZN => n1419);
   U1463 : AOI22_X1 port map( A1 => REGISTERS_0_23_port, A2 => n356, B1 => 
                           REGISTERS_2_23_port, B2 => n319, ZN => n1418);
   U1464 : NAND4_X1 port map( A1 => n1421, A2 => n1420, A3 => n1419, A4 => 
                           n1418, ZN => n1427);
   U1465 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n134_port, B1 
                           => REGISTERS_15_23_port, B2 => n97_port, ZN => n1425
                           );
   U1466 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n208, B1 => 
                           REGISTERS_11_23_port, B2 => n171, ZN => n1424);
   U1467 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n282_port, B1 
                           => REGISTERS_14_23_port, B2 => n245_port, ZN => 
                           n1423);
   U1468 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n356, B1 => 
                           REGISTERS_10_23_port, B2 => n319, ZN => n1422);
   U1469 : NAND4_X1 port map( A1 => n1425, A2 => n1424, A3 => n1423, A4 => 
                           n1422, ZN => n1426);
   U1470 : AOI22_X1 port map( A1 => n1427, A2 => n27, B1 => n1426, B2 => n24, 
                           ZN => n1428);
   U1471 : OAI221_X1 port map( B1 => n2271, B2 => n1430, C1 => n2269, C2 => 
                           n1429, A => n1428, ZN => N136);
   U1472 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n135_port, B1 
                           => REGISTERS_23_24_port, B2 => n98_port, ZN => n1434
                           );
   U1473 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n209, B1 => 
                           REGISTERS_19_24_port, B2 => n172, ZN => n1433);
   U1474 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n283_port, B1 
                           => REGISTERS_22_24_port, B2 => n246_port, ZN => 
                           n1432);
   U1475 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n357, B1 => 
                           REGISTERS_18_24_port, B2 => n320, ZN => n1431);
   U1476 : AND4_X1 port map( A1 => n1434, A2 => n1433, A3 => n1432, A4 => n1431
                           , ZN => n1451);
   U1477 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n135_port, B1 
                           => REGISTERS_31_24_port, B2 => n98_port, ZN => n1438
                           );
   U1478 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n209, B1 => 
                           REGISTERS_27_24_port, B2 => n172, ZN => n1437);
   U1479 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n283_port, B1 
                           => REGISTERS_30_24_port, B2 => n246_port, ZN => 
                           n1436);
   U1480 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n357, B1 => 
                           REGISTERS_26_24_port, B2 => n320, ZN => n1435);
   U1481 : AND4_X1 port map( A1 => n1438, A2 => n1437, A3 => n1436, A4 => n1435
                           , ZN => n1450);
   U1482 : AOI22_X1 port map( A1 => REGISTERS_5_24_port, A2 => n135_port, B1 =>
                           REGISTERS_7_24_port, B2 => n98_port, ZN => n1442);
   U1483 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n209, B1 => 
                           REGISTERS_3_24_port, B2 => n172, ZN => n1441);
   U1484 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n283_port, B1 =>
                           REGISTERS_6_24_port, B2 => n246_port, ZN => n1440);
   U1485 : AOI22_X1 port map( A1 => REGISTERS_0_24_port, A2 => n357, B1 => 
                           REGISTERS_2_24_port, B2 => n320, ZN => n1439);
   U1486 : NAND4_X1 port map( A1 => n1442, A2 => n1441, A3 => n1440, A4 => 
                           n1439, ZN => n1448);
   U1487 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n135_port, B1 
                           => REGISTERS_15_24_port, B2 => n98_port, ZN => n1446
                           );
   U1488 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n209, B1 => 
                           REGISTERS_11_24_port, B2 => n172, ZN => n1445);
   U1489 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n283_port, B1 
                           => REGISTERS_14_24_port, B2 => n246_port, ZN => 
                           n1444);
   U1490 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n357, B1 => 
                           REGISTERS_10_24_port, B2 => n320, ZN => n1443);
   U1491 : NAND4_X1 port map( A1 => n1446, A2 => n1445, A3 => n1444, A4 => 
                           n1443, ZN => n1447);
   U1492 : AOI22_X1 port map( A1 => n1448, A2 => n27, B1 => n1447, B2 => n24, 
                           ZN => n1449);
   U1493 : OAI221_X1 port map( B1 => n2271, B2 => n1451, C1 => n2269, C2 => 
                           n1450, A => n1449, ZN => N135);
   U1494 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n135_port, B1 
                           => REGISTERS_23_25_port, B2 => n98_port, ZN => n1455
                           );
   U1495 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n209, B1 => 
                           REGISTERS_19_25_port, B2 => n172, ZN => n1454);
   U1496 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n283_port, B1 
                           => REGISTERS_22_25_port, B2 => n246_port, ZN => 
                           n1453);
   U1497 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n357, B1 => 
                           REGISTERS_18_25_port, B2 => n320, ZN => n1452);
   U1498 : AND4_X1 port map( A1 => n1455, A2 => n1454, A3 => n1453, A4 => n1452
                           , ZN => n1472);
   U1499 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n135_port, B1 
                           => REGISTERS_31_25_port, B2 => n98_port, ZN => n1459
                           );
   U1500 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n209, B1 => 
                           REGISTERS_27_25_port, B2 => n172, ZN => n1458);
   U1501 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n283_port, B1 
                           => REGISTERS_30_25_port, B2 => n246_port, ZN => 
                           n1457);
   U1502 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n357, B1 => 
                           REGISTERS_26_25_port, B2 => n320, ZN => n1456);
   U1503 : AND4_X1 port map( A1 => n1459, A2 => n1458, A3 => n1457, A4 => n1456
                           , ZN => n1471);
   U1504 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n135_port, B1 =>
                           REGISTERS_7_25_port, B2 => n98_port, ZN => n1463);
   U1505 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n209, B1 => 
                           REGISTERS_3_25_port, B2 => n172, ZN => n1462);
   U1506 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n283_port, B1 =>
                           REGISTERS_6_25_port, B2 => n246_port, ZN => n1461);
   U1507 : AOI22_X1 port map( A1 => REGISTERS_0_25_port, A2 => n357, B1 => 
                           REGISTERS_2_25_port, B2 => n320, ZN => n1460);
   U1508 : NAND4_X1 port map( A1 => n1463, A2 => n1462, A3 => n1461, A4 => 
                           n1460, ZN => n1469);
   U1509 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n135_port, B1 
                           => REGISTERS_15_25_port, B2 => n98_port, ZN => n1467
                           );
   U1510 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n209, B1 => 
                           REGISTERS_11_25_port, B2 => n172, ZN => n1466);
   U1511 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n283_port, B1 
                           => REGISTERS_14_25_port, B2 => n246_port, ZN => 
                           n1465);
   U1512 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n357, B1 => 
                           REGISTERS_10_25_port, B2 => n320, ZN => n1464);
   U1513 : NAND4_X1 port map( A1 => n1467, A2 => n1466, A3 => n1465, A4 => 
                           n1464, ZN => n1468);
   U1514 : AOI22_X1 port map( A1 => n1469, A2 => n27, B1 => n1468, B2 => n24, 
                           ZN => n1470);
   U1515 : OAI221_X1 port map( B1 => n2271, B2 => n1472, C1 => n2269, C2 => 
                           n1471, A => n1470, ZN => N134);
   U1516 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n135_port, B1 
                           => REGISTERS_23_26_port, B2 => n98_port, ZN => n1476
                           );
   U1517 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n209, B1 => 
                           REGISTERS_19_26_port, B2 => n172, ZN => n1475);
   U1518 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n283_port, B1 
                           => REGISTERS_22_26_port, B2 => n246_port, ZN => 
                           n1474);
   U1519 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n357, B1 => 
                           REGISTERS_18_26_port, B2 => n320, ZN => n1473);
   U1520 : AND4_X1 port map( A1 => n1476, A2 => n1475, A3 => n1474, A4 => n1473
                           , ZN => n1493);
   U1521 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n135_port, B1 
                           => REGISTERS_31_26_port, B2 => n98_port, ZN => n1480
                           );
   U1522 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n209, B1 => 
                           REGISTERS_27_26_port, B2 => n172, ZN => n1479);
   U1523 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n283_port, B1 
                           => REGISTERS_30_26_port, B2 => n246_port, ZN => 
                           n1478);
   U1524 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n357, B1 => 
                           REGISTERS_26_26_port, B2 => n320, ZN => n1477);
   U1525 : AND4_X1 port map( A1 => n1480, A2 => n1479, A3 => n1478, A4 => n1477
                           , ZN => n1492);
   U1526 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n135_port, B1 =>
                           REGISTERS_7_26_port, B2 => n98_port, ZN => n1484);
   U1527 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n209, B1 => 
                           REGISTERS_3_26_port, B2 => n172, ZN => n1483);
   U1528 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n283_port, B1 =>
                           REGISTERS_6_26_port, B2 => n246_port, ZN => n1482);
   U1529 : AOI22_X1 port map( A1 => REGISTERS_0_26_port, A2 => n357, B1 => 
                           REGISTERS_2_26_port, B2 => n320, ZN => n1481);
   U1530 : NAND4_X1 port map( A1 => n1484, A2 => n1483, A3 => n1482, A4 => 
                           n1481, ZN => n1490);
   U1531 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n135_port, B1 
                           => REGISTERS_15_26_port, B2 => n98_port, ZN => n1488
                           );
   U1532 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n209, B1 => 
                           REGISTERS_11_26_port, B2 => n172, ZN => n1487);
   U1533 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n283_port, B1 
                           => REGISTERS_14_26_port, B2 => n246_port, ZN => 
                           n1486);
   U1534 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n357, B1 => 
                           REGISTERS_10_26_port, B2 => n320, ZN => n1485);
   U1535 : NAND4_X1 port map( A1 => n1488, A2 => n1487, A3 => n1486, A4 => 
                           n1485, ZN => n1489);
   U1536 : AOI22_X1 port map( A1 => n1490, A2 => n27, B1 => n1489, B2 => n24, 
                           ZN => n1491);
   U1537 : OAI221_X1 port map( B1 => n2271, B2 => n1493, C1 => n2269, C2 => 
                           n1492, A => n1491, ZN => N133);
   U1538 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n136_port, B1 
                           => REGISTERS_23_27_port, B2 => n99_port, ZN => n1497
                           );
   U1539 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n210, B1 => 
                           REGISTERS_19_27_port, B2 => n173, ZN => n1496);
   U1540 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n284_port, B1 
                           => REGISTERS_22_27_port, B2 => n247_port, ZN => 
                           n1495);
   U1541 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n358, B1 => 
                           REGISTERS_18_27_port, B2 => n321, ZN => n1494);
   U1542 : AND4_X1 port map( A1 => n1497, A2 => n1496, A3 => n1495, A4 => n1494
                           , ZN => n1514);
   U1543 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n136_port, B1 
                           => REGISTERS_31_27_port, B2 => n99_port, ZN => n1501
                           );
   U1544 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n210, B1 => 
                           REGISTERS_27_27_port, B2 => n173, ZN => n1500);
   U1545 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n284_port, B1 
                           => REGISTERS_30_27_port, B2 => n247_port, ZN => 
                           n1499);
   U1546 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n358, B1 => 
                           REGISTERS_26_27_port, B2 => n321, ZN => n1498);
   U1547 : AND4_X1 port map( A1 => n1501, A2 => n1500, A3 => n1499, A4 => n1498
                           , ZN => n1513);
   U1548 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n136_port, B1 =>
                           REGISTERS_7_27_port, B2 => n99_port, ZN => n1505);
   U1549 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n210, B1 => 
                           REGISTERS_3_27_port, B2 => n173, ZN => n1504);
   U1550 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n284_port, B1 =>
                           REGISTERS_6_27_port, B2 => n247_port, ZN => n1503);
   U1551 : AOI22_X1 port map( A1 => REGISTERS_0_27_port, A2 => n358, B1 => 
                           REGISTERS_2_27_port, B2 => n321, ZN => n1502);
   U1552 : NAND4_X1 port map( A1 => n1505, A2 => n1504, A3 => n1503, A4 => 
                           n1502, ZN => n1511);
   U1553 : AOI22_X1 port map( A1 => REGISTERS_13_27_port, A2 => n136_port, B1 
                           => REGISTERS_15_27_port, B2 => n99_port, ZN => n1509
                           );
   U1554 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n210, B1 => 
                           REGISTERS_11_27_port, B2 => n173, ZN => n1508);
   U1555 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n284_port, B1 
                           => REGISTERS_14_27_port, B2 => n247_port, ZN => 
                           n1507);
   U1556 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n358, B1 => 
                           REGISTERS_10_27_port, B2 => n321, ZN => n1506);
   U1557 : NAND4_X1 port map( A1 => n1509, A2 => n1508, A3 => n1507, A4 => 
                           n1506, ZN => n1510);
   U1558 : AOI22_X1 port map( A1 => n1511, A2 => n27, B1 => n1510, B2 => n24, 
                           ZN => n1512);
   U1559 : OAI221_X1 port map( B1 => n2271, B2 => n1514, C1 => n2269, C2 => 
                           n1513, A => n1512, ZN => N132);
   U1560 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n136_port, B1 
                           => REGISTERS_23_28_port, B2 => n99_port, ZN => n1518
                           );
   U1561 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n210, B1 => 
                           REGISTERS_19_28_port, B2 => n173, ZN => n1517);
   U1562 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n284_port, B1 
                           => REGISTERS_22_28_port, B2 => n247_port, ZN => 
                           n1516);
   U1563 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n358, B1 => 
                           REGISTERS_18_28_port, B2 => n321, ZN => n1515);
   U1564 : AND4_X1 port map( A1 => n1518, A2 => n1517, A3 => n1516, A4 => n1515
                           , ZN => n1535);
   U1565 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n136_port, B1 
                           => REGISTERS_31_28_port, B2 => n99_port, ZN => n1522
                           );
   U1566 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n210, B1 => 
                           REGISTERS_27_28_port, B2 => n173, ZN => n1521);
   U1567 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n284_port, B1 
                           => REGISTERS_30_28_port, B2 => n247_port, ZN => 
                           n1520);
   U1568 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n358, B1 => 
                           REGISTERS_26_28_port, B2 => n321, ZN => n1519);
   U1569 : AND4_X1 port map( A1 => n1522, A2 => n1521, A3 => n1520, A4 => n1519
                           , ZN => n1534);
   U1570 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n136_port, B1 =>
                           REGISTERS_7_28_port, B2 => n99_port, ZN => n1526);
   U1571 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n210, B1 => 
                           REGISTERS_3_28_port, B2 => n173, ZN => n1525);
   U1572 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n284_port, B1 =>
                           REGISTERS_6_28_port, B2 => n247_port, ZN => n1524);
   U1573 : AOI22_X1 port map( A1 => REGISTERS_0_28_port, A2 => n358, B1 => 
                           REGISTERS_2_28_port, B2 => n321, ZN => n1523);
   U1574 : NAND4_X1 port map( A1 => n1526, A2 => n1525, A3 => n1524, A4 => 
                           n1523, ZN => n1532);
   U1575 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n136_port, B1 
                           => REGISTERS_15_28_port, B2 => n99_port, ZN => n1530
                           );
   U1576 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n210, B1 => 
                           REGISTERS_11_28_port, B2 => n173, ZN => n1529);
   U1577 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n284_port, B1 
                           => REGISTERS_14_28_port, B2 => n247_port, ZN => 
                           n1528);
   U1578 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n358, B1 => 
                           REGISTERS_10_28_port, B2 => n321, ZN => n1527);
   U1579 : NAND4_X1 port map( A1 => n1530, A2 => n1529, A3 => n1528, A4 => 
                           n1527, ZN => n1531);
   U1580 : AOI22_X1 port map( A1 => n1532, A2 => n27, B1 => n1531, B2 => n24, 
                           ZN => n1533);
   U1581 : OAI221_X1 port map( B1 => n2271, B2 => n1535, C1 => n2269, C2 => 
                           n1534, A => n1533, ZN => N131);
   U1582 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n136_port, B1 
                           => REGISTERS_23_29_port, B2 => n99_port, ZN => n1539
                           );
   U1583 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n210, B1 => 
                           REGISTERS_19_29_port, B2 => n173, ZN => n1538);
   U1584 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n284_port, B1 
                           => REGISTERS_22_29_port, B2 => n247_port, ZN => 
                           n1537);
   U1585 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n358, B1 => 
                           REGISTERS_18_29_port, B2 => n321, ZN => n1536);
   U1586 : AND4_X1 port map( A1 => n1539, A2 => n1538, A3 => n1537, A4 => n1536
                           , ZN => n1556);
   U1587 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n136_port, B1 
                           => REGISTERS_31_29_port, B2 => n99_port, ZN => n1543
                           );
   U1588 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n210, B1 => 
                           REGISTERS_27_29_port, B2 => n173, ZN => n1542);
   U1589 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n284_port, B1 
                           => REGISTERS_30_29_port, B2 => n247_port, ZN => 
                           n1541);
   U1590 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n358, B1 => 
                           REGISTERS_26_29_port, B2 => n321, ZN => n1540);
   U1591 : AND4_X1 port map( A1 => n1543, A2 => n1542, A3 => n1541, A4 => n1540
                           , ZN => n1555);
   U1592 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n136_port, B1 =>
                           REGISTERS_7_29_port, B2 => n99_port, ZN => n1547);
   U1593 : AOI22_X1 port map( A1 => REGISTERS_1_29_port, A2 => n210, B1 => 
                           REGISTERS_3_29_port, B2 => n173, ZN => n1546);
   U1594 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n284_port, B1 =>
                           REGISTERS_6_29_port, B2 => n247_port, ZN => n1545);
   U1595 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n358, B1 => 
                           REGISTERS_2_29_port, B2 => n321, ZN => n1544);
   U1596 : NAND4_X1 port map( A1 => n1547, A2 => n1546, A3 => n1545, A4 => 
                           n1544, ZN => n1553);
   U1597 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n136_port, B1 
                           => REGISTERS_15_29_port, B2 => n99_port, ZN => n1551
                           );
   U1598 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n210, B1 => 
                           REGISTERS_11_29_port, B2 => n173, ZN => n1550);
   U1599 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n284_port, B1 
                           => REGISTERS_14_29_port, B2 => n247_port, ZN => 
                           n1549);
   U1600 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n358, B1 => 
                           REGISTERS_10_29_port, B2 => n321, ZN => n1548);
   U1601 : NAND4_X1 port map( A1 => n1551, A2 => n1550, A3 => n1549, A4 => 
                           n1548, ZN => n1552);
   U1602 : AOI22_X1 port map( A1 => n1553, A2 => n27, B1 => n1552, B2 => n24, 
                           ZN => n1554);
   U1603 : OAI221_X1 port map( B1 => n2271, B2 => n1556, C1 => n2269, C2 => 
                           n1555, A => n1554, ZN => N130);
   U1604 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n137_port, B1 
                           => REGISTERS_23_30_port, B2 => n100_port, ZN => 
                           n1560);
   U1605 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n211, B1 => 
                           REGISTERS_19_30_port, B2 => n174, ZN => n1559);
   U1606 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n285_port, B1 
                           => REGISTERS_22_30_port, B2 => n248_port, ZN => 
                           n1558);
   U1607 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n359, B1 => 
                           REGISTERS_18_30_port, B2 => n322, ZN => n1557);
   U1608 : AND4_X1 port map( A1 => n1560, A2 => n1559, A3 => n1558, A4 => n1557
                           , ZN => n1577);
   U1609 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n137_port, B1 
                           => REGISTERS_31_30_port, B2 => n100_port, ZN => 
                           n1564);
   U1610 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n211, B1 => 
                           REGISTERS_27_30_port, B2 => n174, ZN => n1563);
   U1611 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n285_port, B1 
                           => REGISTERS_30_30_port, B2 => n248_port, ZN => 
                           n1562);
   U1612 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n359, B1 => 
                           REGISTERS_26_30_port, B2 => n322, ZN => n1561);
   U1613 : AND4_X1 port map( A1 => n1564, A2 => n1563, A3 => n1562, A4 => n1561
                           , ZN => n1576);
   U1614 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n137_port, B1 =>
                           REGISTERS_7_30_port, B2 => n100_port, ZN => n1568);
   U1615 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n211, B1 => 
                           REGISTERS_3_30_port, B2 => n174, ZN => n1567);
   U1616 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n285_port, B1 =>
                           REGISTERS_6_30_port, B2 => n248_port, ZN => n1566);
   U1617 : AOI22_X1 port map( A1 => REGISTERS_0_30_port, A2 => n359, B1 => 
                           REGISTERS_2_30_port, B2 => n322, ZN => n1565);
   U1618 : NAND4_X1 port map( A1 => n1568, A2 => n1567, A3 => n1566, A4 => 
                           n1565, ZN => n1574);
   U1619 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n137_port, B1 
                           => REGISTERS_15_30_port, B2 => n100_port, ZN => 
                           n1572);
   U1620 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n211, B1 => 
                           REGISTERS_11_30_port, B2 => n174, ZN => n1571);
   U1621 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n285_port, B1 
                           => REGISTERS_14_30_port, B2 => n248_port, ZN => 
                           n1570);
   U1622 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n359, B1 => 
                           REGISTERS_10_30_port, B2 => n322, ZN => n1569);
   U1623 : NAND4_X1 port map( A1 => n1572, A2 => n1571, A3 => n1570, A4 => 
                           n1569, ZN => n1573);
   U1624 : AOI22_X1 port map( A1 => n1574, A2 => n27, B1 => n1573, B2 => n24, 
                           ZN => n1575);
   U1625 : OAI221_X1 port map( B1 => n2271, B2 => n1577, C1 => n2269, C2 => 
                           n1576, A => n1575, ZN => N129);
   U1626 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n137_port, B1 
                           => REGISTERS_23_31_port, B2 => n100_port, ZN => 
                           n1581);
   U1627 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n211, B1 => 
                           REGISTERS_19_31_port, B2 => n174, ZN => n1580);
   U1628 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n285_port, B1 
                           => REGISTERS_22_31_port, B2 => n248_port, ZN => 
                           n1579);
   U1629 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n359, B1 => 
                           REGISTERS_18_31_port, B2 => n322, ZN => n1578);
   U1630 : AND4_X1 port map( A1 => n1581, A2 => n1580, A3 => n1579, A4 => n1578
                           , ZN => n1598);
   U1631 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n137_port, B1 
                           => REGISTERS_31_31_port, B2 => n100_port, ZN => 
                           n1585);
   U1632 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n211, B1 => 
                           REGISTERS_27_31_port, B2 => n174, ZN => n1584);
   U1633 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n285_port, B1 
                           => REGISTERS_30_31_port, B2 => n248_port, ZN => 
                           n1583);
   U1634 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n359, B1 => 
                           REGISTERS_26_31_port, B2 => n322, ZN => n1582);
   U1635 : AND4_X1 port map( A1 => n1585, A2 => n1584, A3 => n1583, A4 => n1582
                           , ZN => n1597);
   U1636 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n137_port, B1 =>
                           REGISTERS_7_31_port, B2 => n100_port, ZN => n1589);
   U1637 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n211, B1 => 
                           REGISTERS_3_31_port, B2 => n174, ZN => n1588);
   U1638 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n285_port, B1 =>
                           REGISTERS_6_31_port, B2 => n248_port, ZN => n1587);
   U1639 : AOI22_X1 port map( A1 => REGISTERS_0_31_port, A2 => n359, B1 => 
                           REGISTERS_2_31_port, B2 => n322, ZN => n1586);
   U1640 : NAND4_X1 port map( A1 => n1589, A2 => n1588, A3 => n1587, A4 => 
                           n1586, ZN => n1595);
   U1641 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n137_port, B1 
                           => REGISTERS_15_31_port, B2 => n100_port, ZN => 
                           n1593);
   U1642 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n211, B1 => 
                           REGISTERS_11_31_port, B2 => n174, ZN => n1592);
   U1643 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n285_port, B1 
                           => REGISTERS_14_31_port, B2 => n248_port, ZN => 
                           n1591);
   U1644 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n359, B1 => 
                           REGISTERS_10_31_port, B2 => n322, ZN => n1590);
   U1645 : NAND4_X1 port map( A1 => n1593, A2 => n1592, A3 => n1591, A4 => 
                           n1590, ZN => n1594);
   U1646 : AOI22_X1 port map( A1 => n1595, A2 => n27, B1 => n1594, B2 => n24, 
                           ZN => n1596);
   U1647 : OAI221_X1 port map( B1 => n2271, B2 => n1598, C1 => n2269, C2 => 
                           n1597, A => n1596, ZN => N128);
   U1648 : AOI22_X1 port map( A1 => REGISTERS_21_32_port, A2 => n137_port, B1 
                           => REGISTERS_23_32_port, B2 => n100_port, ZN => 
                           n1602);
   U1649 : AOI22_X1 port map( A1 => REGISTERS_17_32_port, A2 => n211, B1 => 
                           REGISTERS_19_32_port, B2 => n174, ZN => n1601);
   U1650 : AOI22_X1 port map( A1 => REGISTERS_20_32_port, A2 => n285_port, B1 
                           => REGISTERS_22_32_port, B2 => n248_port, ZN => 
                           n1600);
   U1651 : AOI22_X1 port map( A1 => REGISTERS_16_32_port, A2 => n359, B1 => 
                           REGISTERS_18_32_port, B2 => n322, ZN => n1599);
   U1652 : AND4_X1 port map( A1 => n1602, A2 => n1601, A3 => n1600, A4 => n1599
                           , ZN => n1619);
   U1653 : AOI22_X1 port map( A1 => REGISTERS_29_32_port, A2 => n137_port, B1 
                           => REGISTERS_31_32_port, B2 => n100_port, ZN => 
                           n1606);
   U1654 : AOI22_X1 port map( A1 => REGISTERS_25_32_port, A2 => n211, B1 => 
                           REGISTERS_27_32_port, B2 => n174, ZN => n1605);
   U1655 : AOI22_X1 port map( A1 => REGISTERS_28_32_port, A2 => n285_port, B1 
                           => REGISTERS_30_32_port, B2 => n248_port, ZN => 
                           n1604);
   U1656 : AOI22_X1 port map( A1 => REGISTERS_24_32_port, A2 => n359, B1 => 
                           REGISTERS_26_32_port, B2 => n322, ZN => n1603);
   U1657 : AND4_X1 port map( A1 => n1606, A2 => n1605, A3 => n1604, A4 => n1603
                           , ZN => n1618);
   U1658 : AOI22_X1 port map( A1 => REGISTERS_5_32_port, A2 => n137_port, B1 =>
                           REGISTERS_7_32_port, B2 => n100_port, ZN => n1610);
   U1659 : AOI22_X1 port map( A1 => REGISTERS_1_32_port, A2 => n211, B1 => 
                           REGISTERS_3_32_port, B2 => n174, ZN => n1609);
   U1660 : AOI22_X1 port map( A1 => REGISTERS_4_32_port, A2 => n285_port, B1 =>
                           REGISTERS_6_32_port, B2 => n248_port, ZN => n1608);
   U1661 : AOI22_X1 port map( A1 => REGISTERS_0_32_port, A2 => n359, B1 => 
                           REGISTERS_2_32_port, B2 => n322, ZN => n1607);
   U1662 : NAND4_X1 port map( A1 => n1610, A2 => n1609, A3 => n1608, A4 => 
                           n1607, ZN => n1616);
   U1663 : AOI22_X1 port map( A1 => REGISTERS_13_32_port, A2 => n137_port, B1 
                           => REGISTERS_15_32_port, B2 => n100_port, ZN => 
                           n1614);
   U1664 : AOI22_X1 port map( A1 => REGISTERS_9_32_port, A2 => n211, B1 => 
                           REGISTERS_11_32_port, B2 => n174, ZN => n1613);
   U1665 : AOI22_X1 port map( A1 => REGISTERS_12_32_port, A2 => n285_port, B1 
                           => REGISTERS_14_32_port, B2 => n248_port, ZN => 
                           n1612);
   U1666 : AOI22_X1 port map( A1 => REGISTERS_8_32_port, A2 => n359, B1 => 
                           REGISTERS_10_32_port, B2 => n322, ZN => n1611);
   U1667 : NAND4_X1 port map( A1 => n1614, A2 => n1613, A3 => n1612, A4 => 
                           n1611, ZN => n1615);
   U1668 : AOI22_X1 port map( A1 => n1616, A2 => n27, B1 => n1615, B2 => n24, 
                           ZN => n1617);
   U1669 : OAI221_X1 port map( B1 => n2271, B2 => n1619, C1 => n2269, C2 => 
                           n1618, A => n1617, ZN => N127);
   U1670 : AOI22_X1 port map( A1 => REGISTERS_21_33_port, A2 => n138_port, B1 
                           => REGISTERS_23_33_port, B2 => n101_port, ZN => 
                           n1623);
   U1671 : AOI22_X1 port map( A1 => REGISTERS_17_33_port, A2 => n212, B1 => 
                           REGISTERS_19_33_port, B2 => n175, ZN => n1622);
   U1672 : AOI22_X1 port map( A1 => REGISTERS_20_33_port, A2 => n286_port, B1 
                           => REGISTERS_22_33_port, B2 => n249_port, ZN => 
                           n1621);
   U1673 : AOI22_X1 port map( A1 => REGISTERS_16_33_port, A2 => n360, B1 => 
                           REGISTERS_18_33_port, B2 => n323, ZN => n1620);
   U1674 : AND4_X1 port map( A1 => n1623, A2 => n1622, A3 => n1621, A4 => n1620
                           , ZN => n1640);
   U1675 : AOI22_X1 port map( A1 => REGISTERS_29_33_port, A2 => n138_port, B1 
                           => REGISTERS_31_33_port, B2 => n101_port, ZN => 
                           n1627);
   U1676 : AOI22_X1 port map( A1 => REGISTERS_25_33_port, A2 => n212, B1 => 
                           REGISTERS_27_33_port, B2 => n175, ZN => n1626);
   U1677 : AOI22_X1 port map( A1 => REGISTERS_28_33_port, A2 => n286_port, B1 
                           => REGISTERS_30_33_port, B2 => n249_port, ZN => 
                           n1625);
   U1678 : AOI22_X1 port map( A1 => REGISTERS_24_33_port, A2 => n360, B1 => 
                           REGISTERS_26_33_port, B2 => n323, ZN => n1624);
   U1679 : AND4_X1 port map( A1 => n1627, A2 => n1626, A3 => n1625, A4 => n1624
                           , ZN => n1639);
   U1680 : AOI22_X1 port map( A1 => REGISTERS_5_33_port, A2 => n138_port, B1 =>
                           REGISTERS_7_33_port, B2 => n101_port, ZN => n1631);
   U1681 : AOI22_X1 port map( A1 => REGISTERS_1_33_port, A2 => n212, B1 => 
                           REGISTERS_3_33_port, B2 => n175, ZN => n1630);
   U1682 : AOI22_X1 port map( A1 => REGISTERS_4_33_port, A2 => n286_port, B1 =>
                           REGISTERS_6_33_port, B2 => n249_port, ZN => n1629);
   U1683 : AOI22_X1 port map( A1 => REGISTERS_0_33_port, A2 => n360, B1 => 
                           REGISTERS_2_33_port, B2 => n323, ZN => n1628);
   U1684 : NAND4_X1 port map( A1 => n1631, A2 => n1630, A3 => n1629, A4 => 
                           n1628, ZN => n1637);
   U1685 : AOI22_X1 port map( A1 => REGISTERS_13_33_port, A2 => n138_port, B1 
                           => REGISTERS_15_33_port, B2 => n101_port, ZN => 
                           n1635);
   U1686 : AOI22_X1 port map( A1 => REGISTERS_9_33_port, A2 => n212, B1 => 
                           REGISTERS_11_33_port, B2 => n175, ZN => n1634);
   U1687 : AOI22_X1 port map( A1 => REGISTERS_12_33_port, A2 => n286_port, B1 
                           => REGISTERS_14_33_port, B2 => n249_port, ZN => 
                           n1633);
   U1688 : AOI22_X1 port map( A1 => REGISTERS_8_33_port, A2 => n360, B1 => 
                           REGISTERS_10_33_port, B2 => n323, ZN => n1632);
   U1689 : NAND4_X1 port map( A1 => n1635, A2 => n1634, A3 => n1633, A4 => 
                           n1632, ZN => n1636);
   U1690 : AOI22_X1 port map( A1 => n1637, A2 => n27, B1 => n1636, B2 => n24, 
                           ZN => n1638);
   U1691 : OAI221_X1 port map( B1 => n2271, B2 => n1640, C1 => n2269, C2 => 
                           n1639, A => n1638, ZN => N126);
   U1692 : AOI22_X1 port map( A1 => REGISTERS_21_34_port, A2 => n138_port, B1 
                           => REGISTERS_23_34_port, B2 => n101_port, ZN => 
                           n1644);
   U1693 : AOI22_X1 port map( A1 => REGISTERS_17_34_port, A2 => n212, B1 => 
                           REGISTERS_19_34_port, B2 => n175, ZN => n1643);
   U1694 : AOI22_X1 port map( A1 => REGISTERS_20_34_port, A2 => n286_port, B1 
                           => REGISTERS_22_34_port, B2 => n249_port, ZN => 
                           n1642);
   U1695 : AOI22_X1 port map( A1 => REGISTERS_16_34_port, A2 => n360, B1 => 
                           REGISTERS_18_34_port, B2 => n323, ZN => n1641);
   U1696 : AND4_X1 port map( A1 => n1644, A2 => n1643, A3 => n1642, A4 => n1641
                           , ZN => n1661);
   U1697 : AOI22_X1 port map( A1 => REGISTERS_29_34_port, A2 => n138_port, B1 
                           => REGISTERS_31_34_port, B2 => n101_port, ZN => 
                           n1648);
   U1698 : AOI22_X1 port map( A1 => REGISTERS_25_34_port, A2 => n212, B1 => 
                           REGISTERS_27_34_port, B2 => n175, ZN => n1647);
   U1699 : AOI22_X1 port map( A1 => REGISTERS_28_34_port, A2 => n286_port, B1 
                           => REGISTERS_30_34_port, B2 => n249_port, ZN => 
                           n1646);
   U1700 : AOI22_X1 port map( A1 => REGISTERS_24_34_port, A2 => n360, B1 => 
                           REGISTERS_26_34_port, B2 => n323, ZN => n1645);
   U1701 : AND4_X1 port map( A1 => n1648, A2 => n1647, A3 => n1646, A4 => n1645
                           , ZN => n1660);
   U1702 : AOI22_X1 port map( A1 => REGISTERS_5_34_port, A2 => n138_port, B1 =>
                           REGISTERS_7_34_port, B2 => n101_port, ZN => n1652);
   U1703 : AOI22_X1 port map( A1 => REGISTERS_1_34_port, A2 => n212, B1 => 
                           REGISTERS_3_34_port, B2 => n175, ZN => n1651);
   U1704 : AOI22_X1 port map( A1 => REGISTERS_4_34_port, A2 => n286_port, B1 =>
                           REGISTERS_6_34_port, B2 => n249_port, ZN => n1650);
   U1705 : AOI22_X1 port map( A1 => REGISTERS_0_34_port, A2 => n360, B1 => 
                           REGISTERS_2_34_port, B2 => n323, ZN => n1649);
   U1706 : NAND4_X1 port map( A1 => n1652, A2 => n1651, A3 => n1650, A4 => 
                           n1649, ZN => n1658);
   U1707 : AOI22_X1 port map( A1 => REGISTERS_13_34_port, A2 => n138_port, B1 
                           => REGISTERS_15_34_port, B2 => n101_port, ZN => 
                           n1656);
   U1708 : AOI22_X1 port map( A1 => REGISTERS_9_34_port, A2 => n212, B1 => 
                           REGISTERS_11_34_port, B2 => n175, ZN => n1655);
   U1709 : AOI22_X1 port map( A1 => REGISTERS_12_34_port, A2 => n286_port, B1 
                           => REGISTERS_14_34_port, B2 => n249_port, ZN => 
                           n1654);
   U1710 : AOI22_X1 port map( A1 => REGISTERS_8_34_port, A2 => n360, B1 => 
                           REGISTERS_10_34_port, B2 => n323, ZN => n1653);
   U1711 : NAND4_X1 port map( A1 => n1656, A2 => n1655, A3 => n1654, A4 => 
                           n1653, ZN => n1657);
   U1712 : AOI22_X1 port map( A1 => n1658, A2 => n27, B1 => n1657, B2 => n24, 
                           ZN => n1659);
   U1713 : OAI221_X1 port map( B1 => n2271, B2 => n1661, C1 => n2269, C2 => 
                           n1660, A => n1659, ZN => N125);
   U1714 : AOI22_X1 port map( A1 => REGISTERS_21_35_port, A2 => n138_port, B1 
                           => REGISTERS_23_35_port, B2 => n101_port, ZN => 
                           n1665);
   U1715 : AOI22_X1 port map( A1 => REGISTERS_17_35_port, A2 => n212, B1 => 
                           REGISTERS_19_35_port, B2 => n175, ZN => n1664);
   U1716 : AOI22_X1 port map( A1 => REGISTERS_20_35_port, A2 => n286_port, B1 
                           => REGISTERS_22_35_port, B2 => n249_port, ZN => 
                           n1663);
   U1717 : AOI22_X1 port map( A1 => REGISTERS_16_35_port, A2 => n360, B1 => 
                           REGISTERS_18_35_port, B2 => n323, ZN => n1662);
   U1718 : AND4_X1 port map( A1 => n1665, A2 => n1664, A3 => n1663, A4 => n1662
                           , ZN => n1682);
   U1719 : AOI22_X1 port map( A1 => REGISTERS_29_35_port, A2 => n138_port, B1 
                           => REGISTERS_31_35_port, B2 => n101_port, ZN => 
                           n1669);
   U1720 : AOI22_X1 port map( A1 => REGISTERS_25_35_port, A2 => n212, B1 => 
                           REGISTERS_27_35_port, B2 => n175, ZN => n1668);
   U1721 : AOI22_X1 port map( A1 => REGISTERS_28_35_port, A2 => n286_port, B1 
                           => REGISTERS_30_35_port, B2 => n249_port, ZN => 
                           n1667);
   U1722 : AOI22_X1 port map( A1 => REGISTERS_24_35_port, A2 => n360, B1 => 
                           REGISTERS_26_35_port, B2 => n323, ZN => n1666);
   U1723 : AND4_X1 port map( A1 => n1669, A2 => n1668, A3 => n1667, A4 => n1666
                           , ZN => n1681);
   U1724 : AOI22_X1 port map( A1 => REGISTERS_5_35_port, A2 => n138_port, B1 =>
                           REGISTERS_7_35_port, B2 => n101_port, ZN => n1673);
   U1725 : AOI22_X1 port map( A1 => REGISTERS_1_35_port, A2 => n212, B1 => 
                           REGISTERS_3_35_port, B2 => n175, ZN => n1672);
   U1726 : AOI22_X1 port map( A1 => REGISTERS_4_35_port, A2 => n286_port, B1 =>
                           REGISTERS_6_35_port, B2 => n249_port, ZN => n1671);
   U1727 : AOI22_X1 port map( A1 => REGISTERS_0_35_port, A2 => n360, B1 => 
                           REGISTERS_2_35_port, B2 => n323, ZN => n1670);
   U1728 : NAND4_X1 port map( A1 => n1673, A2 => n1672, A3 => n1671, A4 => 
                           n1670, ZN => n1679);
   U1729 : AOI22_X1 port map( A1 => REGISTERS_13_35_port, A2 => n138_port, B1 
                           => REGISTERS_15_35_port, B2 => n101_port, ZN => 
                           n1677);
   U1730 : AOI22_X1 port map( A1 => REGISTERS_9_35_port, A2 => n212, B1 => 
                           REGISTERS_11_35_port, B2 => n175, ZN => n1676);
   U1731 : AOI22_X1 port map( A1 => REGISTERS_12_35_port, A2 => n286_port, B1 
                           => REGISTERS_14_35_port, B2 => n249_port, ZN => 
                           n1675);
   U1732 : AOI22_X1 port map( A1 => REGISTERS_8_35_port, A2 => n360, B1 => 
                           REGISTERS_10_35_port, B2 => n323, ZN => n1674);
   U1733 : NAND4_X1 port map( A1 => n1677, A2 => n1676, A3 => n1675, A4 => 
                           n1674, ZN => n1678);
   U1734 : AOI22_X1 port map( A1 => n1679, A2 => n27, B1 => n1678, B2 => n24, 
                           ZN => n1680);
   U1735 : OAI221_X1 port map( B1 => n2271, B2 => n1682, C1 => n2269, C2 => 
                           n1681, A => n1680, ZN => N124);
   U1736 : AOI22_X1 port map( A1 => REGISTERS_21_36_port, A2 => n139_port, B1 
                           => REGISTERS_23_36_port, B2 => n102_port, ZN => 
                           n1686);
   U1737 : AOI22_X1 port map( A1 => REGISTERS_17_36_port, A2 => n213, B1 => 
                           REGISTERS_19_36_port, B2 => n176, ZN => n1685);
   U1738 : AOI22_X1 port map( A1 => REGISTERS_20_36_port, A2 => n287_port, B1 
                           => REGISTERS_22_36_port, B2 => n250_port, ZN => 
                           n1684);
   U1739 : AOI22_X1 port map( A1 => REGISTERS_16_36_port, A2 => n361, B1 => 
                           REGISTERS_18_36_port, B2 => n324, ZN => n1683);
   U1740 : AND4_X1 port map( A1 => n1686, A2 => n1685, A3 => n1684, A4 => n1683
                           , ZN => n1703);
   U1741 : AOI22_X1 port map( A1 => REGISTERS_29_36_port, A2 => n139_port, B1 
                           => REGISTERS_31_36_port, B2 => n102_port, ZN => 
                           n1690);
   U1742 : AOI22_X1 port map( A1 => REGISTERS_25_36_port, A2 => n213, B1 => 
                           REGISTERS_27_36_port, B2 => n176, ZN => n1689);
   U1743 : AOI22_X1 port map( A1 => REGISTERS_28_36_port, A2 => n287_port, B1 
                           => REGISTERS_30_36_port, B2 => n250_port, ZN => 
                           n1688);
   U1744 : AOI22_X1 port map( A1 => REGISTERS_24_36_port, A2 => n361, B1 => 
                           REGISTERS_26_36_port, B2 => n324, ZN => n1687);
   U1745 : AND4_X1 port map( A1 => n1690, A2 => n1689, A3 => n1688, A4 => n1687
                           , ZN => n1702);
   U1746 : AOI22_X1 port map( A1 => REGISTERS_5_36_port, A2 => n139_port, B1 =>
                           REGISTERS_7_36_port, B2 => n102_port, ZN => n1694);
   U1747 : AOI22_X1 port map( A1 => REGISTERS_1_36_port, A2 => n213, B1 => 
                           REGISTERS_3_36_port, B2 => n176, ZN => n1693);
   U1748 : AOI22_X1 port map( A1 => REGISTERS_4_36_port, A2 => n287_port, B1 =>
                           REGISTERS_6_36_port, B2 => n250_port, ZN => n1692);
   U1749 : AOI22_X1 port map( A1 => REGISTERS_0_36_port, A2 => n361, B1 => 
                           REGISTERS_2_36_port, B2 => n324, ZN => n1691);
   U1750 : NAND4_X1 port map( A1 => n1694, A2 => n1693, A3 => n1692, A4 => 
                           n1691, ZN => n1700);
   U1751 : AOI22_X1 port map( A1 => REGISTERS_13_36_port, A2 => n139_port, B1 
                           => REGISTERS_15_36_port, B2 => n102_port, ZN => 
                           n1698);
   U1752 : AOI22_X1 port map( A1 => REGISTERS_9_36_port, A2 => n213, B1 => 
                           REGISTERS_11_36_port, B2 => n176, ZN => n1697);
   U1753 : AOI22_X1 port map( A1 => REGISTERS_12_36_port, A2 => n287_port, B1 
                           => REGISTERS_14_36_port, B2 => n250_port, ZN => 
                           n1696);
   U1754 : AOI22_X1 port map( A1 => REGISTERS_8_36_port, A2 => n361, B1 => 
                           REGISTERS_10_36_port, B2 => n324, ZN => n1695);
   U1755 : NAND4_X1 port map( A1 => n1698, A2 => n1697, A3 => n1696, A4 => 
                           n1695, ZN => n1699);
   U1756 : AOI22_X1 port map( A1 => n1700, A2 => n27, B1 => n1699, B2 => n24, 
                           ZN => n1701);
   U1757 : OAI221_X1 port map( B1 => n2271, B2 => n1703, C1 => n2269, C2 => 
                           n1702, A => n1701, ZN => N123);
   U1758 : AOI22_X1 port map( A1 => REGISTERS_21_37_port, A2 => n139_port, B1 
                           => REGISTERS_23_37_port, B2 => n102_port, ZN => 
                           n1707);
   U1759 : AOI22_X1 port map( A1 => REGISTERS_17_37_port, A2 => n213, B1 => 
                           REGISTERS_19_37_port, B2 => n176, ZN => n1706);
   U1760 : AOI22_X1 port map( A1 => REGISTERS_20_37_port, A2 => n287_port, B1 
                           => REGISTERS_22_37_port, B2 => n250_port, ZN => 
                           n1705);
   U1761 : AOI22_X1 port map( A1 => REGISTERS_16_37_port, A2 => n361, B1 => 
                           REGISTERS_18_37_port, B2 => n324, ZN => n1704);
   U1762 : AND4_X1 port map( A1 => n1707, A2 => n1706, A3 => n1705, A4 => n1704
                           , ZN => n1724);
   U1763 : AOI22_X1 port map( A1 => REGISTERS_29_37_port, A2 => n139_port, B1 
                           => REGISTERS_31_37_port, B2 => n102_port, ZN => 
                           n1711);
   U1764 : AOI22_X1 port map( A1 => REGISTERS_25_37_port, A2 => n213, B1 => 
                           REGISTERS_27_37_port, B2 => n176, ZN => n1710);
   U1765 : AOI22_X1 port map( A1 => REGISTERS_28_37_port, A2 => n287_port, B1 
                           => REGISTERS_30_37_port, B2 => n250_port, ZN => 
                           n1709);
   U1766 : AOI22_X1 port map( A1 => REGISTERS_24_37_port, A2 => n361, B1 => 
                           REGISTERS_26_37_port, B2 => n324, ZN => n1708);
   U1767 : AND4_X1 port map( A1 => n1711, A2 => n1710, A3 => n1709, A4 => n1708
                           , ZN => n1723);
   U1768 : AOI22_X1 port map( A1 => REGISTERS_5_37_port, A2 => n139_port, B1 =>
                           REGISTERS_7_37_port, B2 => n102_port, ZN => n1715);
   U1769 : AOI22_X1 port map( A1 => REGISTERS_1_37_port, A2 => n213, B1 => 
                           REGISTERS_3_37_port, B2 => n176, ZN => n1714);
   U1770 : AOI22_X1 port map( A1 => REGISTERS_4_37_port, A2 => n287_port, B1 =>
                           REGISTERS_6_37_port, B2 => n250_port, ZN => n1713);
   U1771 : AOI22_X1 port map( A1 => REGISTERS_0_37_port, A2 => n361, B1 => 
                           REGISTERS_2_37_port, B2 => n324, ZN => n1712);
   U1772 : NAND4_X1 port map( A1 => n1715, A2 => n1714, A3 => n1713, A4 => 
                           n1712, ZN => n1721);
   U1773 : AOI22_X1 port map( A1 => REGISTERS_13_37_port, A2 => n139_port, B1 
                           => REGISTERS_15_37_port, B2 => n102_port, ZN => 
                           n1719);
   U1774 : AOI22_X1 port map( A1 => REGISTERS_9_37_port, A2 => n213, B1 => 
                           REGISTERS_11_37_port, B2 => n176, ZN => n1718);
   U1775 : AOI22_X1 port map( A1 => REGISTERS_12_37_port, A2 => n287_port, B1 
                           => REGISTERS_14_37_port, B2 => n250_port, ZN => 
                           n1717);
   U1776 : AOI22_X1 port map( A1 => REGISTERS_8_37_port, A2 => n361, B1 => 
                           REGISTERS_10_37_port, B2 => n324, ZN => n1716);
   U1777 : NAND4_X1 port map( A1 => n1719, A2 => n1718, A3 => n1717, A4 => 
                           n1716, ZN => n1720);
   U1778 : AOI22_X1 port map( A1 => n1721, A2 => n27, B1 => n1720, B2 => n24, 
                           ZN => n1722);
   U1779 : OAI221_X1 port map( B1 => n2271, B2 => n1724, C1 => n2269, C2 => 
                           n1723, A => n1722, ZN => N122);
   U1780 : AOI22_X1 port map( A1 => REGISTERS_21_38_port, A2 => n139_port, B1 
                           => REGISTERS_23_38_port, B2 => n102_port, ZN => 
                           n1728);
   U1781 : AOI22_X1 port map( A1 => REGISTERS_17_38_port, A2 => n213, B1 => 
                           REGISTERS_19_38_port, B2 => n176, ZN => n1727);
   U1782 : AOI22_X1 port map( A1 => REGISTERS_20_38_port, A2 => n287_port, B1 
                           => REGISTERS_22_38_port, B2 => n250_port, ZN => 
                           n1726);
   U1783 : AOI22_X1 port map( A1 => REGISTERS_16_38_port, A2 => n361, B1 => 
                           REGISTERS_18_38_port, B2 => n324, ZN => n1725);
   U1784 : AND4_X1 port map( A1 => n1728, A2 => n1727, A3 => n1726, A4 => n1725
                           , ZN => n1745);
   U1785 : AOI22_X1 port map( A1 => REGISTERS_29_38_port, A2 => n139_port, B1 
                           => REGISTERS_31_38_port, B2 => n102_port, ZN => 
                           n1732);
   U1786 : AOI22_X1 port map( A1 => REGISTERS_25_38_port, A2 => n213, B1 => 
                           REGISTERS_27_38_port, B2 => n176, ZN => n1731);
   U1787 : AOI22_X1 port map( A1 => REGISTERS_28_38_port, A2 => n287_port, B1 
                           => REGISTERS_30_38_port, B2 => n250_port, ZN => 
                           n1730);
   U1788 : AOI22_X1 port map( A1 => REGISTERS_24_38_port, A2 => n361, B1 => 
                           REGISTERS_26_38_port, B2 => n324, ZN => n1729);
   U1789 : AND4_X1 port map( A1 => n1732, A2 => n1731, A3 => n1730, A4 => n1729
                           , ZN => n1744);
   U1790 : AOI22_X1 port map( A1 => REGISTERS_5_38_port, A2 => n139_port, B1 =>
                           REGISTERS_7_38_port, B2 => n102_port, ZN => n1736);
   U1791 : AOI22_X1 port map( A1 => REGISTERS_1_38_port, A2 => n213, B1 => 
                           REGISTERS_3_38_port, B2 => n176, ZN => n1735);
   U1792 : AOI22_X1 port map( A1 => REGISTERS_4_38_port, A2 => n287_port, B1 =>
                           REGISTERS_6_38_port, B2 => n250_port, ZN => n1734);
   U1793 : AOI22_X1 port map( A1 => REGISTERS_0_38_port, A2 => n361, B1 => 
                           REGISTERS_2_38_port, B2 => n324, ZN => n1733);
   U1794 : NAND4_X1 port map( A1 => n1736, A2 => n1735, A3 => n1734, A4 => 
                           n1733, ZN => n1742);
   U1795 : AOI22_X1 port map( A1 => REGISTERS_13_38_port, A2 => n139_port, B1 
                           => REGISTERS_15_38_port, B2 => n102_port, ZN => 
                           n1740);
   U1796 : AOI22_X1 port map( A1 => REGISTERS_9_38_port, A2 => n213, B1 => 
                           REGISTERS_11_38_port, B2 => n176, ZN => n1739);
   U1797 : AOI22_X1 port map( A1 => REGISTERS_12_38_port, A2 => n287_port, B1 
                           => REGISTERS_14_38_port, B2 => n250_port, ZN => 
                           n1738);
   U1798 : AOI22_X1 port map( A1 => REGISTERS_8_38_port, A2 => n361, B1 => 
                           REGISTERS_10_38_port, B2 => n324, ZN => n1737);
   U1799 : NAND4_X1 port map( A1 => n1740, A2 => n1739, A3 => n1738, A4 => 
                           n1737, ZN => n1741);
   U1800 : AOI22_X1 port map( A1 => n1742, A2 => n27, B1 => n1741, B2 => n24, 
                           ZN => n1743);
   U1801 : OAI221_X1 port map( B1 => n2271, B2 => n1745, C1 => n2269, C2 => 
                           n1744, A => n1743, ZN => N121);
   U1802 : AOI22_X1 port map( A1 => REGISTERS_21_39_port, A2 => n140_port, B1 
                           => REGISTERS_23_39_port, B2 => n103_port, ZN => 
                           n1749);
   U1803 : AOI22_X1 port map( A1 => REGISTERS_17_39_port, A2 => n214, B1 => 
                           REGISTERS_19_39_port, B2 => n177, ZN => n1748);
   U1804 : AOI22_X1 port map( A1 => REGISTERS_20_39_port, A2 => n288_port, B1 
                           => REGISTERS_22_39_port, B2 => n251_port, ZN => 
                           n1747);
   U1805 : AOI22_X1 port map( A1 => REGISTERS_16_39_port, A2 => n362, B1 => 
                           REGISTERS_18_39_port, B2 => n325, ZN => n1746);
   U1806 : AND4_X1 port map( A1 => n1749, A2 => n1748, A3 => n1747, A4 => n1746
                           , ZN => n1766);
   U1807 : AOI22_X1 port map( A1 => REGISTERS_29_39_port, A2 => n140_port, B1 
                           => REGISTERS_31_39_port, B2 => n103_port, ZN => 
                           n1753);
   U1808 : AOI22_X1 port map( A1 => REGISTERS_25_39_port, A2 => n214, B1 => 
                           REGISTERS_27_39_port, B2 => n177, ZN => n1752);
   U1809 : AOI22_X1 port map( A1 => REGISTERS_28_39_port, A2 => n288_port, B1 
                           => REGISTERS_30_39_port, B2 => n251_port, ZN => 
                           n1751);
   U1810 : AOI22_X1 port map( A1 => REGISTERS_24_39_port, A2 => n362, B1 => 
                           REGISTERS_26_39_port, B2 => n325, ZN => n1750);
   U1811 : AND4_X1 port map( A1 => n1753, A2 => n1752, A3 => n1751, A4 => n1750
                           , ZN => n1765);
   U1812 : AOI22_X1 port map( A1 => REGISTERS_5_39_port, A2 => n140_port, B1 =>
                           REGISTERS_7_39_port, B2 => n103_port, ZN => n1757);
   U1813 : AOI22_X1 port map( A1 => REGISTERS_1_39_port, A2 => n214, B1 => 
                           REGISTERS_3_39_port, B2 => n177, ZN => n1756);
   U1814 : AOI22_X1 port map( A1 => REGISTERS_4_39_port, A2 => n288_port, B1 =>
                           REGISTERS_6_39_port, B2 => n251_port, ZN => n1755);
   U1815 : AOI22_X1 port map( A1 => REGISTERS_0_39_port, A2 => n362, B1 => 
                           REGISTERS_2_39_port, B2 => n325, ZN => n1754);
   U1816 : NAND4_X1 port map( A1 => n1757, A2 => n1756, A3 => n1755, A4 => 
                           n1754, ZN => n1763);
   U1817 : AOI22_X1 port map( A1 => REGISTERS_13_39_port, A2 => n140_port, B1 
                           => REGISTERS_15_39_port, B2 => n103_port, ZN => 
                           n1761);
   U1818 : AOI22_X1 port map( A1 => REGISTERS_9_39_port, A2 => n214, B1 => 
                           REGISTERS_11_39_port, B2 => n177, ZN => n1760);
   U1819 : AOI22_X1 port map( A1 => REGISTERS_12_39_port, A2 => n288_port, B1 
                           => REGISTERS_14_39_port, B2 => n251_port, ZN => 
                           n1759);
   U1820 : AOI22_X1 port map( A1 => REGISTERS_8_39_port, A2 => n362, B1 => 
                           REGISTERS_10_39_port, B2 => n325, ZN => n1758);
   U1821 : NAND4_X1 port map( A1 => n1761, A2 => n1760, A3 => n1759, A4 => 
                           n1758, ZN => n1762);
   U1822 : AOI22_X1 port map( A1 => n1763, A2 => n27, B1 => n1762, B2 => n24, 
                           ZN => n1764);
   U1823 : OAI221_X1 port map( B1 => n2271, B2 => n1766, C1 => n2269, C2 => 
                           n1765, A => n1764, ZN => N120);
   U1824 : AOI22_X1 port map( A1 => REGISTERS_21_40_port, A2 => n140_port, B1 
                           => REGISTERS_23_40_port, B2 => n103_port, ZN => 
                           n1770);
   U1825 : AOI22_X1 port map( A1 => REGISTERS_17_40_port, A2 => n214, B1 => 
                           REGISTERS_19_40_port, B2 => n177, ZN => n1769);
   U1826 : AOI22_X1 port map( A1 => REGISTERS_20_40_port, A2 => n288_port, B1 
                           => REGISTERS_22_40_port, B2 => n251_port, ZN => 
                           n1768);
   U1827 : AOI22_X1 port map( A1 => REGISTERS_16_40_port, A2 => n362, B1 => 
                           REGISTERS_18_40_port, B2 => n325, ZN => n1767);
   U1828 : AND4_X1 port map( A1 => n1770, A2 => n1769, A3 => n1768, A4 => n1767
                           , ZN => n1787);
   U1829 : AOI22_X1 port map( A1 => REGISTERS_29_40_port, A2 => n140_port, B1 
                           => REGISTERS_31_40_port, B2 => n103_port, ZN => 
                           n1774);
   U1830 : AOI22_X1 port map( A1 => REGISTERS_25_40_port, A2 => n214, B1 => 
                           REGISTERS_27_40_port, B2 => n177, ZN => n1773);
   U1831 : AOI22_X1 port map( A1 => REGISTERS_28_40_port, A2 => n288_port, B1 
                           => REGISTERS_30_40_port, B2 => n251_port, ZN => 
                           n1772);
   U1832 : AOI22_X1 port map( A1 => REGISTERS_24_40_port, A2 => n362, B1 => 
                           REGISTERS_26_40_port, B2 => n325, ZN => n1771);
   U1833 : AND4_X1 port map( A1 => n1774, A2 => n1773, A3 => n1772, A4 => n1771
                           , ZN => n1786);
   U1834 : AOI22_X1 port map( A1 => REGISTERS_5_40_port, A2 => n140_port, B1 =>
                           REGISTERS_7_40_port, B2 => n103_port, ZN => n1778);
   U1835 : AOI22_X1 port map( A1 => REGISTERS_1_40_port, A2 => n214, B1 => 
                           REGISTERS_3_40_port, B2 => n177, ZN => n1777);
   U1836 : AOI22_X1 port map( A1 => REGISTERS_4_40_port, A2 => n288_port, B1 =>
                           REGISTERS_6_40_port, B2 => n251_port, ZN => n1776);
   U1837 : AOI22_X1 port map( A1 => REGISTERS_0_40_port, A2 => n362, B1 => 
                           REGISTERS_2_40_port, B2 => n325, ZN => n1775);
   U1838 : NAND4_X1 port map( A1 => n1778, A2 => n1777, A3 => n1776, A4 => 
                           n1775, ZN => n1784);
   U1839 : AOI22_X1 port map( A1 => REGISTERS_13_40_port, A2 => n140_port, B1 
                           => REGISTERS_15_40_port, B2 => n103_port, ZN => 
                           n1782);
   U1840 : AOI22_X1 port map( A1 => REGISTERS_9_40_port, A2 => n214, B1 => 
                           REGISTERS_11_40_port, B2 => n177, ZN => n1781);
   U1841 : AOI22_X1 port map( A1 => REGISTERS_12_40_port, A2 => n288_port, B1 
                           => REGISTERS_14_40_port, B2 => n251_port, ZN => 
                           n1780);
   U1842 : AOI22_X1 port map( A1 => REGISTERS_8_40_port, A2 => n362, B1 => 
                           REGISTERS_10_40_port, B2 => n325, ZN => n1779);
   U1843 : NAND4_X1 port map( A1 => n1782, A2 => n1781, A3 => n1780, A4 => 
                           n1779, ZN => n1783);
   U1844 : AOI22_X1 port map( A1 => n1784, A2 => n27, B1 => n1783, B2 => n24, 
                           ZN => n1785);
   U1845 : OAI221_X1 port map( B1 => n2271, B2 => n1787, C1 => n2269, C2 => 
                           n1786, A => n1785, ZN => N119);
   U1846 : AOI22_X1 port map( A1 => REGISTERS_21_41_port, A2 => n140_port, B1 
                           => REGISTERS_23_41_port, B2 => n103_port, ZN => 
                           n1791);
   U1847 : AOI22_X1 port map( A1 => REGISTERS_17_41_port, A2 => n214, B1 => 
                           REGISTERS_19_41_port, B2 => n177, ZN => n1790);
   U1848 : AOI22_X1 port map( A1 => REGISTERS_20_41_port, A2 => n288_port, B1 
                           => REGISTERS_22_41_port, B2 => n251_port, ZN => 
                           n1789);
   U1849 : AOI22_X1 port map( A1 => REGISTERS_16_41_port, A2 => n362, B1 => 
                           REGISTERS_18_41_port, B2 => n325, ZN => n1788);
   U1850 : AND4_X1 port map( A1 => n1791, A2 => n1790, A3 => n1789, A4 => n1788
                           , ZN => n1808);
   U1851 : AOI22_X1 port map( A1 => REGISTERS_29_41_port, A2 => n140_port, B1 
                           => REGISTERS_31_41_port, B2 => n103_port, ZN => 
                           n1795);
   U1852 : AOI22_X1 port map( A1 => REGISTERS_25_41_port, A2 => n214, B1 => 
                           REGISTERS_27_41_port, B2 => n177, ZN => n1794);
   U1853 : AOI22_X1 port map( A1 => REGISTERS_28_41_port, A2 => n288_port, B1 
                           => REGISTERS_30_41_port, B2 => n251_port, ZN => 
                           n1793);
   U1854 : AOI22_X1 port map( A1 => REGISTERS_24_41_port, A2 => n362, B1 => 
                           REGISTERS_26_41_port, B2 => n325, ZN => n1792);
   U1855 : AND4_X1 port map( A1 => n1795, A2 => n1794, A3 => n1793, A4 => n1792
                           , ZN => n1807);
   U1856 : AOI22_X1 port map( A1 => REGISTERS_5_41_port, A2 => n140_port, B1 =>
                           REGISTERS_7_41_port, B2 => n103_port, ZN => n1799);
   U1857 : AOI22_X1 port map( A1 => REGISTERS_1_41_port, A2 => n214, B1 => 
                           REGISTERS_3_41_port, B2 => n177, ZN => n1798);
   U1858 : AOI22_X1 port map( A1 => REGISTERS_4_41_port, A2 => n288_port, B1 =>
                           REGISTERS_6_41_port, B2 => n251_port, ZN => n1797);
   U1859 : AOI22_X1 port map( A1 => REGISTERS_0_41_port, A2 => n362, B1 => 
                           REGISTERS_2_41_port, B2 => n325, ZN => n1796);
   U1860 : NAND4_X1 port map( A1 => n1799, A2 => n1798, A3 => n1797, A4 => 
                           n1796, ZN => n1805);
   U1861 : AOI22_X1 port map( A1 => REGISTERS_13_41_port, A2 => n140_port, B1 
                           => REGISTERS_15_41_port, B2 => n103_port, ZN => 
                           n1803);
   U1862 : AOI22_X1 port map( A1 => REGISTERS_9_41_port, A2 => n214, B1 => 
                           REGISTERS_11_41_port, B2 => n177, ZN => n1802);
   U1863 : AOI22_X1 port map( A1 => REGISTERS_12_41_port, A2 => n288_port, B1 
                           => REGISTERS_14_41_port, B2 => n251_port, ZN => 
                           n1801);
   U1864 : AOI22_X1 port map( A1 => REGISTERS_8_41_port, A2 => n362, B1 => 
                           REGISTERS_10_41_port, B2 => n325, ZN => n1800);
   U1865 : NAND4_X1 port map( A1 => n1803, A2 => n1802, A3 => n1801, A4 => 
                           n1800, ZN => n1804);
   U1866 : AOI22_X1 port map( A1 => n1805, A2 => n27, B1 => n1804, B2 => n24, 
                           ZN => n1806);
   U1867 : OAI221_X1 port map( B1 => n2271, B2 => n1808, C1 => n2269, C2 => 
                           n1807, A => n1806, ZN => N118);
   U1868 : AOI22_X1 port map( A1 => REGISTERS_21_42_port, A2 => n141_port, B1 
                           => REGISTERS_23_42_port, B2 => n104_port, ZN => 
                           n1812);
   U1869 : AOI22_X1 port map( A1 => REGISTERS_17_42_port, A2 => n215, B1 => 
                           REGISTERS_19_42_port, B2 => n178, ZN => n1811);
   U1870 : AOI22_X1 port map( A1 => REGISTERS_20_42_port, A2 => n289, B1 => 
                           REGISTERS_22_42_port, B2 => n252_port, ZN => n1810);
   U1871 : AOI22_X1 port map( A1 => REGISTERS_16_42_port, A2 => n363, B1 => 
                           REGISTERS_18_42_port, B2 => n326, ZN => n1809);
   U1872 : AND4_X1 port map( A1 => n1812, A2 => n1811, A3 => n1810, A4 => n1809
                           , ZN => n1829);
   U1873 : AOI22_X1 port map( A1 => REGISTERS_29_42_port, A2 => n141_port, B1 
                           => REGISTERS_31_42_port, B2 => n104_port, ZN => 
                           n1816);
   U1874 : AOI22_X1 port map( A1 => REGISTERS_25_42_port, A2 => n215, B1 => 
                           REGISTERS_27_42_port, B2 => n178, ZN => n1815);
   U1875 : AOI22_X1 port map( A1 => REGISTERS_28_42_port, A2 => n289, B1 => 
                           REGISTERS_30_42_port, B2 => n252_port, ZN => n1814);
   U1876 : AOI22_X1 port map( A1 => REGISTERS_24_42_port, A2 => n363, B1 => 
                           REGISTERS_26_42_port, B2 => n326, ZN => n1813);
   U1877 : AND4_X1 port map( A1 => n1816, A2 => n1815, A3 => n1814, A4 => n1813
                           , ZN => n1828);
   U1878 : AOI22_X1 port map( A1 => REGISTERS_5_42_port, A2 => n141_port, B1 =>
                           REGISTERS_7_42_port, B2 => n104_port, ZN => n1820);
   U1879 : AOI22_X1 port map( A1 => REGISTERS_1_42_port, A2 => n215, B1 => 
                           REGISTERS_3_42_port, B2 => n178, ZN => n1819);
   U1880 : AOI22_X1 port map( A1 => REGISTERS_4_42_port, A2 => n289, B1 => 
                           REGISTERS_6_42_port, B2 => n252_port, ZN => n1818);
   U1881 : AOI22_X1 port map( A1 => REGISTERS_0_42_port, A2 => n363, B1 => 
                           REGISTERS_2_42_port, B2 => n326, ZN => n1817);
   U1882 : NAND4_X1 port map( A1 => n1820, A2 => n1819, A3 => n1818, A4 => 
                           n1817, ZN => n1826);
   U1883 : AOI22_X1 port map( A1 => REGISTERS_13_42_port, A2 => n141_port, B1 
                           => REGISTERS_15_42_port, B2 => n104_port, ZN => 
                           n1824);
   U1884 : AOI22_X1 port map( A1 => REGISTERS_9_42_port, A2 => n215, B1 => 
                           REGISTERS_11_42_port, B2 => n178, ZN => n1823);
   U1885 : AOI22_X1 port map( A1 => REGISTERS_12_42_port, A2 => n289, B1 => 
                           REGISTERS_14_42_port, B2 => n252_port, ZN => n1822);
   U1886 : AOI22_X1 port map( A1 => REGISTERS_8_42_port, A2 => n363, B1 => 
                           REGISTERS_10_42_port, B2 => n326, ZN => n1821);
   U1887 : NAND4_X1 port map( A1 => n1824, A2 => n1823, A3 => n1822, A4 => 
                           n1821, ZN => n1825);
   U1888 : AOI22_X1 port map( A1 => n1826, A2 => n27, B1 => n1825, B2 => n24, 
                           ZN => n1827);
   U1889 : OAI221_X1 port map( B1 => n2271, B2 => n1829, C1 => n2269, C2 => 
                           n1828, A => n1827, ZN => N117);
   U1890 : AOI22_X1 port map( A1 => REGISTERS_21_43_port, A2 => n141_port, B1 
                           => REGISTERS_23_43_port, B2 => n104_port, ZN => 
                           n1833);
   U1891 : AOI22_X1 port map( A1 => REGISTERS_17_43_port, A2 => n215, B1 => 
                           REGISTERS_19_43_port, B2 => n178, ZN => n1832);
   U1892 : AOI22_X1 port map( A1 => REGISTERS_20_43_port, A2 => n289, B1 => 
                           REGISTERS_22_43_port, B2 => n252_port, ZN => n1831);
   U1893 : AOI22_X1 port map( A1 => REGISTERS_16_43_port, A2 => n363, B1 => 
                           REGISTERS_18_43_port, B2 => n326, ZN => n1830);
   U1894 : AND4_X1 port map( A1 => n1833, A2 => n1832, A3 => n1831, A4 => n1830
                           , ZN => n1850);
   U1895 : AOI22_X1 port map( A1 => REGISTERS_29_43_port, A2 => n141_port, B1 
                           => REGISTERS_31_43_port, B2 => n104_port, ZN => 
                           n1837);
   U1896 : AOI22_X1 port map( A1 => REGISTERS_25_43_port, A2 => n215, B1 => 
                           REGISTERS_27_43_port, B2 => n178, ZN => n1836);
   U1897 : AOI22_X1 port map( A1 => REGISTERS_28_43_port, A2 => n289, B1 => 
                           REGISTERS_30_43_port, B2 => n252_port, ZN => n1835);
   U1898 : AOI22_X1 port map( A1 => REGISTERS_24_43_port, A2 => n363, B1 => 
                           REGISTERS_26_43_port, B2 => n326, ZN => n1834);
   U1899 : AND4_X1 port map( A1 => n1837, A2 => n1836, A3 => n1835, A4 => n1834
                           , ZN => n1849);
   U1900 : AOI22_X1 port map( A1 => REGISTERS_5_43_port, A2 => n141_port, B1 =>
                           REGISTERS_7_43_port, B2 => n104_port, ZN => n1841);
   U1901 : AOI22_X1 port map( A1 => REGISTERS_1_43_port, A2 => n215, B1 => 
                           REGISTERS_3_43_port, B2 => n178, ZN => n1840);
   U1902 : AOI22_X1 port map( A1 => REGISTERS_4_43_port, A2 => n289, B1 => 
                           REGISTERS_6_43_port, B2 => n252_port, ZN => n1839);
   U1903 : AOI22_X1 port map( A1 => REGISTERS_0_43_port, A2 => n363, B1 => 
                           REGISTERS_2_43_port, B2 => n326, ZN => n1838);
   U1904 : NAND4_X1 port map( A1 => n1841, A2 => n1840, A3 => n1839, A4 => 
                           n1838, ZN => n1847);
   U1905 : AOI22_X1 port map( A1 => REGISTERS_13_43_port, A2 => n141_port, B1 
                           => REGISTERS_15_43_port, B2 => n104_port, ZN => 
                           n1845);
   U1906 : AOI22_X1 port map( A1 => REGISTERS_9_43_port, A2 => n215, B1 => 
                           REGISTERS_11_43_port, B2 => n178, ZN => n1844);
   U1907 : AOI22_X1 port map( A1 => REGISTERS_12_43_port, A2 => n289, B1 => 
                           REGISTERS_14_43_port, B2 => n252_port, ZN => n1843);
   U1908 : AOI22_X1 port map( A1 => REGISTERS_8_43_port, A2 => n363, B1 => 
                           REGISTERS_10_43_port, B2 => n326, ZN => n1842);
   U1909 : NAND4_X1 port map( A1 => n1845, A2 => n1844, A3 => n1843, A4 => 
                           n1842, ZN => n1846);
   U1910 : AOI22_X1 port map( A1 => n1847, A2 => n27, B1 => n1846, B2 => n24, 
                           ZN => n1848);
   U1911 : OAI221_X1 port map( B1 => n2271, B2 => n1850, C1 => n2269, C2 => 
                           n1849, A => n1848, ZN => N116);
   U1912 : AOI22_X1 port map( A1 => REGISTERS_21_44_port, A2 => n141_port, B1 
                           => REGISTERS_23_44_port, B2 => n104_port, ZN => 
                           n1854);
   U1913 : AOI22_X1 port map( A1 => REGISTERS_17_44_port, A2 => n215, B1 => 
                           REGISTERS_19_44_port, B2 => n178, ZN => n1853);
   U1914 : AOI22_X1 port map( A1 => REGISTERS_20_44_port, A2 => n289, B1 => 
                           REGISTERS_22_44_port, B2 => n252_port, ZN => n1852);
   U1915 : AOI22_X1 port map( A1 => REGISTERS_16_44_port, A2 => n363, B1 => 
                           REGISTERS_18_44_port, B2 => n326, ZN => n1851);
   U1916 : AND4_X1 port map( A1 => n1854, A2 => n1853, A3 => n1852, A4 => n1851
                           , ZN => n1871);
   U1917 : AOI22_X1 port map( A1 => REGISTERS_29_44_port, A2 => n141_port, B1 
                           => REGISTERS_31_44_port, B2 => n104_port, ZN => 
                           n1858);
   U1918 : AOI22_X1 port map( A1 => REGISTERS_25_44_port, A2 => n215, B1 => 
                           REGISTERS_27_44_port, B2 => n178, ZN => n1857);
   U1919 : AOI22_X1 port map( A1 => REGISTERS_28_44_port, A2 => n289, B1 => 
                           REGISTERS_30_44_port, B2 => n252_port, ZN => n1856);
   U1920 : AOI22_X1 port map( A1 => REGISTERS_24_44_port, A2 => n363, B1 => 
                           REGISTERS_26_44_port, B2 => n326, ZN => n1855);
   U1921 : AND4_X1 port map( A1 => n1858, A2 => n1857, A3 => n1856, A4 => n1855
                           , ZN => n1870);
   U1922 : AOI22_X1 port map( A1 => REGISTERS_5_44_port, A2 => n141_port, B1 =>
                           REGISTERS_7_44_port, B2 => n104_port, ZN => n1862);
   U1923 : AOI22_X1 port map( A1 => REGISTERS_1_44_port, A2 => n215, B1 => 
                           REGISTERS_3_44_port, B2 => n178, ZN => n1861);
   U1924 : AOI22_X1 port map( A1 => REGISTERS_4_44_port, A2 => n289, B1 => 
                           REGISTERS_6_44_port, B2 => n252_port, ZN => n1860);
   U1925 : AOI22_X1 port map( A1 => REGISTERS_0_44_port, A2 => n363, B1 => 
                           REGISTERS_2_44_port, B2 => n326, ZN => n1859);
   U1926 : NAND4_X1 port map( A1 => n1862, A2 => n1861, A3 => n1860, A4 => 
                           n1859, ZN => n1868);
   U1927 : AOI22_X1 port map( A1 => REGISTERS_13_44_port, A2 => n141_port, B1 
                           => REGISTERS_15_44_port, B2 => n104_port, ZN => 
                           n1866);
   U1928 : AOI22_X1 port map( A1 => REGISTERS_9_44_port, A2 => n215, B1 => 
                           REGISTERS_11_44_port, B2 => n178, ZN => n1865);
   U1929 : AOI22_X1 port map( A1 => REGISTERS_12_44_port, A2 => n289, B1 => 
                           REGISTERS_14_44_port, B2 => n252_port, ZN => n1864);
   U1930 : AOI22_X1 port map( A1 => REGISTERS_8_44_port, A2 => n363, B1 => 
                           REGISTERS_10_44_port, B2 => n326, ZN => n1863);
   U1931 : NAND4_X1 port map( A1 => n1866, A2 => n1865, A3 => n1864, A4 => 
                           n1863, ZN => n1867);
   U1932 : AOI22_X1 port map( A1 => n1868, A2 => n27, B1 => n1867, B2 => n24, 
                           ZN => n1869);
   U1933 : OAI221_X1 port map( B1 => n2271, B2 => n1871, C1 => n2269, C2 => 
                           n1870, A => n1869, ZN => N115);
   U1934 : AOI22_X1 port map( A1 => REGISTERS_21_45_port, A2 => n142_port, B1 
                           => REGISTERS_23_45_port, B2 => n105_port, ZN => 
                           n1875);
   U1935 : AOI22_X1 port map( A1 => REGISTERS_17_45_port, A2 => n216, B1 => 
                           REGISTERS_19_45_port, B2 => n179, ZN => n1874);
   U1936 : AOI22_X1 port map( A1 => REGISTERS_20_45_port, A2 => n290, B1 => 
                           REGISTERS_22_45_port, B2 => n253_port, ZN => n1873);
   U1937 : AOI22_X1 port map( A1 => REGISTERS_16_45_port, A2 => n364, B1 => 
                           REGISTERS_18_45_port, B2 => n327, ZN => n1872);
   U1938 : AND4_X1 port map( A1 => n1875, A2 => n1874, A3 => n1873, A4 => n1872
                           , ZN => n1892);
   U1939 : AOI22_X1 port map( A1 => REGISTERS_29_45_port, A2 => n142_port, B1 
                           => REGISTERS_31_45_port, B2 => n105_port, ZN => 
                           n1879);
   U1940 : AOI22_X1 port map( A1 => REGISTERS_25_45_port, A2 => n216, B1 => 
                           REGISTERS_27_45_port, B2 => n179, ZN => n1878);
   U1941 : AOI22_X1 port map( A1 => REGISTERS_28_45_port, A2 => n290, B1 => 
                           REGISTERS_30_45_port, B2 => n253_port, ZN => n1877);
   U1942 : AOI22_X1 port map( A1 => REGISTERS_24_45_port, A2 => n364, B1 => 
                           REGISTERS_26_45_port, B2 => n327, ZN => n1876);
   U1943 : AND4_X1 port map( A1 => n1879, A2 => n1878, A3 => n1877, A4 => n1876
                           , ZN => n1891);
   U1944 : AOI22_X1 port map( A1 => REGISTERS_5_45_port, A2 => n142_port, B1 =>
                           REGISTERS_7_45_port, B2 => n105_port, ZN => n1883);
   U1945 : AOI22_X1 port map( A1 => REGISTERS_1_45_port, A2 => n216, B1 => 
                           REGISTERS_3_45_port, B2 => n179, ZN => n1882);
   U1946 : AOI22_X1 port map( A1 => REGISTERS_4_45_port, A2 => n290, B1 => 
                           REGISTERS_6_45_port, B2 => n253_port, ZN => n1881);
   U1947 : AOI22_X1 port map( A1 => REGISTERS_0_45_port, A2 => n364, B1 => 
                           REGISTERS_2_45_port, B2 => n327, ZN => n1880);
   U1948 : NAND4_X1 port map( A1 => n1883, A2 => n1882, A3 => n1881, A4 => 
                           n1880, ZN => n1889);
   U1949 : AOI22_X1 port map( A1 => REGISTERS_13_45_port, A2 => n142_port, B1 
                           => REGISTERS_15_45_port, B2 => n105_port, ZN => 
                           n1887);
   U1950 : AOI22_X1 port map( A1 => REGISTERS_9_45_port, A2 => n216, B1 => 
                           REGISTERS_11_45_port, B2 => n179, ZN => n1886);
   U1951 : AOI22_X1 port map( A1 => REGISTERS_12_45_port, A2 => n290, B1 => 
                           REGISTERS_14_45_port, B2 => n253_port, ZN => n1885);
   U1952 : AOI22_X1 port map( A1 => REGISTERS_8_45_port, A2 => n364, B1 => 
                           REGISTERS_10_45_port, B2 => n327, ZN => n1884);
   U1953 : NAND4_X1 port map( A1 => n1887, A2 => n1886, A3 => n1885, A4 => 
                           n1884, ZN => n1888);
   U1954 : AOI22_X1 port map( A1 => n1889, A2 => n27, B1 => n1888, B2 => n24, 
                           ZN => n1890);
   U1955 : OAI221_X1 port map( B1 => n2271, B2 => n1892, C1 => n2269, C2 => 
                           n1891, A => n1890, ZN => N114);
   U1956 : AOI22_X1 port map( A1 => REGISTERS_21_46_port, A2 => n142_port, B1 
                           => REGISTERS_23_46_port, B2 => n105_port, ZN => 
                           n1896);
   U1957 : AOI22_X1 port map( A1 => REGISTERS_17_46_port, A2 => n216, B1 => 
                           REGISTERS_19_46_port, B2 => n179, ZN => n1895);
   U1958 : AOI22_X1 port map( A1 => REGISTERS_20_46_port, A2 => n290, B1 => 
                           REGISTERS_22_46_port, B2 => n253_port, ZN => n1894);
   U1959 : AOI22_X1 port map( A1 => REGISTERS_16_46_port, A2 => n364, B1 => 
                           REGISTERS_18_46_port, B2 => n327, ZN => n1893);
   U1960 : AND4_X1 port map( A1 => n1896, A2 => n1895, A3 => n1894, A4 => n1893
                           , ZN => n1913);
   U1961 : AOI22_X1 port map( A1 => REGISTERS_29_46_port, A2 => n142_port, B1 
                           => REGISTERS_31_46_port, B2 => n105_port, ZN => 
                           n1900);
   U1962 : AOI22_X1 port map( A1 => REGISTERS_25_46_port, A2 => n216, B1 => 
                           REGISTERS_27_46_port, B2 => n179, ZN => n1899);
   U1963 : AOI22_X1 port map( A1 => REGISTERS_28_46_port, A2 => n290, B1 => 
                           REGISTERS_30_46_port, B2 => n253_port, ZN => n1898);
   U1964 : AOI22_X1 port map( A1 => REGISTERS_24_46_port, A2 => n364, B1 => 
                           REGISTERS_26_46_port, B2 => n327, ZN => n1897);
   U1965 : AND4_X1 port map( A1 => n1900, A2 => n1899, A3 => n1898, A4 => n1897
                           , ZN => n1912);
   U1966 : AOI22_X1 port map( A1 => REGISTERS_5_46_port, A2 => n142_port, B1 =>
                           REGISTERS_7_46_port, B2 => n105_port, ZN => n1904);
   U1967 : AOI22_X1 port map( A1 => REGISTERS_1_46_port, A2 => n216, B1 => 
                           REGISTERS_3_46_port, B2 => n179, ZN => n1903);
   U1968 : AOI22_X1 port map( A1 => REGISTERS_4_46_port, A2 => n290, B1 => 
                           REGISTERS_6_46_port, B2 => n253_port, ZN => n1902);
   U1969 : AOI22_X1 port map( A1 => REGISTERS_0_46_port, A2 => n364, B1 => 
                           REGISTERS_2_46_port, B2 => n327, ZN => n1901);
   U1970 : NAND4_X1 port map( A1 => n1904, A2 => n1903, A3 => n1902, A4 => 
                           n1901, ZN => n1910);
   U1971 : AOI22_X1 port map( A1 => REGISTERS_13_46_port, A2 => n142_port, B1 
                           => REGISTERS_15_46_port, B2 => n105_port, ZN => 
                           n1908);
   U1972 : AOI22_X1 port map( A1 => REGISTERS_9_46_port, A2 => n216, B1 => 
                           REGISTERS_11_46_port, B2 => n179, ZN => n1907);
   U1973 : AOI22_X1 port map( A1 => REGISTERS_12_46_port, A2 => n290, B1 => 
                           REGISTERS_14_46_port, B2 => n253_port, ZN => n1906);
   U1974 : AOI22_X1 port map( A1 => REGISTERS_8_46_port, A2 => n364, B1 => 
                           REGISTERS_10_46_port, B2 => n327, ZN => n1905);
   U1975 : NAND4_X1 port map( A1 => n1908, A2 => n1907, A3 => n1906, A4 => 
                           n1905, ZN => n1909);
   U1976 : AOI22_X1 port map( A1 => n1910, A2 => n27, B1 => n1909, B2 => n24, 
                           ZN => n1911);
   U1977 : OAI221_X1 port map( B1 => n2271, B2 => n1913, C1 => n2269, C2 => 
                           n1912, A => n1911, ZN => N113);
   U1978 : AOI22_X1 port map( A1 => REGISTERS_21_47_port, A2 => n142_port, B1 
                           => REGISTERS_23_47_port, B2 => n105_port, ZN => 
                           n1917);
   U1979 : AOI22_X1 port map( A1 => REGISTERS_17_47_port, A2 => n216, B1 => 
                           REGISTERS_19_47_port, B2 => n179, ZN => n1916);
   U1980 : AOI22_X1 port map( A1 => REGISTERS_20_47_port, A2 => n290, B1 => 
                           REGISTERS_22_47_port, B2 => n253_port, ZN => n1915);
   U1981 : AOI22_X1 port map( A1 => REGISTERS_16_47_port, A2 => n364, B1 => 
                           REGISTERS_18_47_port, B2 => n327, ZN => n1914);
   U1982 : AND4_X1 port map( A1 => n1917, A2 => n1916, A3 => n1915, A4 => n1914
                           , ZN => n1934);
   U1983 : AOI22_X1 port map( A1 => REGISTERS_29_47_port, A2 => n142_port, B1 
                           => REGISTERS_31_47_port, B2 => n105_port, ZN => 
                           n1921);
   U1984 : AOI22_X1 port map( A1 => REGISTERS_25_47_port, A2 => n216, B1 => 
                           REGISTERS_27_47_port, B2 => n179, ZN => n1920);
   U1985 : AOI22_X1 port map( A1 => REGISTERS_28_47_port, A2 => n290, B1 => 
                           REGISTERS_30_47_port, B2 => n253_port, ZN => n1919);
   U1986 : AOI22_X1 port map( A1 => REGISTERS_24_47_port, A2 => n364, B1 => 
                           REGISTERS_26_47_port, B2 => n327, ZN => n1918);
   U1987 : AND4_X1 port map( A1 => n1921, A2 => n1920, A3 => n1919, A4 => n1918
                           , ZN => n1933);
   U1988 : AOI22_X1 port map( A1 => REGISTERS_5_47_port, A2 => n142_port, B1 =>
                           REGISTERS_7_47_port, B2 => n105_port, ZN => n1925);
   U1989 : AOI22_X1 port map( A1 => REGISTERS_1_47_port, A2 => n216, B1 => 
                           REGISTERS_3_47_port, B2 => n179, ZN => n1924);
   U1990 : AOI22_X1 port map( A1 => REGISTERS_4_47_port, A2 => n290, B1 => 
                           REGISTERS_6_47_port, B2 => n253_port, ZN => n1923);
   U1991 : AOI22_X1 port map( A1 => REGISTERS_0_47_port, A2 => n364, B1 => 
                           REGISTERS_2_47_port, B2 => n327, ZN => n1922);
   U1992 : NAND4_X1 port map( A1 => n1925, A2 => n1924, A3 => n1923, A4 => 
                           n1922, ZN => n1931);
   U1993 : AOI22_X1 port map( A1 => REGISTERS_13_47_port, A2 => n142_port, B1 
                           => REGISTERS_15_47_port, B2 => n105_port, ZN => 
                           n1929);
   U1994 : AOI22_X1 port map( A1 => REGISTERS_9_47_port, A2 => n216, B1 => 
                           REGISTERS_11_47_port, B2 => n179, ZN => n1928);
   U1995 : AOI22_X1 port map( A1 => REGISTERS_12_47_port, A2 => n290, B1 => 
                           REGISTERS_14_47_port, B2 => n253_port, ZN => n1927);
   U1996 : AOI22_X1 port map( A1 => REGISTERS_8_47_port, A2 => n364, B1 => 
                           REGISTERS_10_47_port, B2 => n327, ZN => n1926);
   U1997 : NAND4_X1 port map( A1 => n1929, A2 => n1928, A3 => n1927, A4 => 
                           n1926, ZN => n1930);
   U1998 : AOI22_X1 port map( A1 => n1931, A2 => n27, B1 => n1930, B2 => n24, 
                           ZN => n1932);
   U1999 : OAI221_X1 port map( B1 => n2271, B2 => n1934, C1 => n2269, C2 => 
                           n1933, A => n1932, ZN => N112);
   U2000 : AOI22_X1 port map( A1 => REGISTERS_21_48_port, A2 => n143_port, B1 
                           => REGISTERS_23_48_port, B2 => n106_port, ZN => 
                           n1938);
   U2001 : AOI22_X1 port map( A1 => REGISTERS_17_48_port, A2 => n217, B1 => 
                           REGISTERS_19_48_port, B2 => n180, ZN => n1937);
   U2002 : AOI22_X1 port map( A1 => REGISTERS_20_48_port, A2 => n291, B1 => 
                           REGISTERS_22_48_port, B2 => n254_port, ZN => n1936);
   U2003 : AOI22_X1 port map( A1 => REGISTERS_16_48_port, A2 => n365, B1 => 
                           REGISTERS_18_48_port, B2 => n328, ZN => n1935);
   U2004 : AND4_X1 port map( A1 => n1938, A2 => n1937, A3 => n1936, A4 => n1935
                           , ZN => n1955);
   U2005 : AOI22_X1 port map( A1 => REGISTERS_29_48_port, A2 => n143_port, B1 
                           => REGISTERS_31_48_port, B2 => n106_port, ZN => 
                           n1942);
   U2006 : AOI22_X1 port map( A1 => REGISTERS_25_48_port, A2 => n217, B1 => 
                           REGISTERS_27_48_port, B2 => n180, ZN => n1941);
   U2007 : AOI22_X1 port map( A1 => REGISTERS_28_48_port, A2 => n291, B1 => 
                           REGISTERS_30_48_port, B2 => n254_port, ZN => n1940);
   U2008 : AOI22_X1 port map( A1 => REGISTERS_24_48_port, A2 => n365, B1 => 
                           REGISTERS_26_48_port, B2 => n328, ZN => n1939);
   U2009 : AND4_X1 port map( A1 => n1942, A2 => n1941, A3 => n1940, A4 => n1939
                           , ZN => n1954);
   U2010 : AOI22_X1 port map( A1 => REGISTERS_5_48_port, A2 => n143_port, B1 =>
                           REGISTERS_7_48_port, B2 => n106_port, ZN => n1946);
   U2011 : AOI22_X1 port map( A1 => REGISTERS_1_48_port, A2 => n217, B1 => 
                           REGISTERS_3_48_port, B2 => n180, ZN => n1945);
   U2012 : AOI22_X1 port map( A1 => REGISTERS_4_48_port, A2 => n291, B1 => 
                           REGISTERS_6_48_port, B2 => n254_port, ZN => n1944);
   U2013 : AOI22_X1 port map( A1 => REGISTERS_0_48_port, A2 => n365, B1 => 
                           REGISTERS_2_48_port, B2 => n328, ZN => n1943);
   U2014 : NAND4_X1 port map( A1 => n1946, A2 => n1945, A3 => n1944, A4 => 
                           n1943, ZN => n1952);
   U2015 : AOI22_X1 port map( A1 => REGISTERS_13_48_port, A2 => n143_port, B1 
                           => REGISTERS_15_48_port, B2 => n106_port, ZN => 
                           n1950);
   U2016 : AOI22_X1 port map( A1 => REGISTERS_9_48_port, A2 => n217, B1 => 
                           REGISTERS_11_48_port, B2 => n180, ZN => n1949);
   U2017 : AOI22_X1 port map( A1 => REGISTERS_12_48_port, A2 => n291, B1 => 
                           REGISTERS_14_48_port, B2 => n254_port, ZN => n1948);
   U2018 : AOI22_X1 port map( A1 => REGISTERS_8_48_port, A2 => n365, B1 => 
                           REGISTERS_10_48_port, B2 => n328, ZN => n1947);
   U2019 : NAND4_X1 port map( A1 => n1950, A2 => n1949, A3 => n1948, A4 => 
                           n1947, ZN => n1951);
   U2020 : AOI22_X1 port map( A1 => n1952, A2 => n27, B1 => n1951, B2 => n24, 
                           ZN => n1953);
   U2021 : OAI221_X1 port map( B1 => n2271, B2 => n1955, C1 => n2269, C2 => 
                           n1954, A => n1953, ZN => N111);
   U2022 : AOI22_X1 port map( A1 => REGISTERS_21_49_port, A2 => n143_port, B1 
                           => REGISTERS_23_49_port, B2 => n106_port, ZN => 
                           n1959);
   U2023 : AOI22_X1 port map( A1 => REGISTERS_17_49_port, A2 => n217, B1 => 
                           REGISTERS_19_49_port, B2 => n180, ZN => n1958);
   U2024 : AOI22_X1 port map( A1 => REGISTERS_20_49_port, A2 => n291, B1 => 
                           REGISTERS_22_49_port, B2 => n254_port, ZN => n1957);
   U2025 : AOI22_X1 port map( A1 => REGISTERS_16_49_port, A2 => n365, B1 => 
                           REGISTERS_18_49_port, B2 => n328, ZN => n1956);
   U2026 : AND4_X1 port map( A1 => n1959, A2 => n1958, A3 => n1957, A4 => n1956
                           , ZN => n1976);
   U2027 : AOI22_X1 port map( A1 => REGISTERS_29_49_port, A2 => n143_port, B1 
                           => REGISTERS_31_49_port, B2 => n106_port, ZN => 
                           n1963);
   U2028 : AOI22_X1 port map( A1 => REGISTERS_25_49_port, A2 => n217, B1 => 
                           REGISTERS_27_49_port, B2 => n180, ZN => n1962);
   U2029 : AOI22_X1 port map( A1 => REGISTERS_28_49_port, A2 => n291, B1 => 
                           REGISTERS_30_49_port, B2 => n254_port, ZN => n1961);
   U2030 : AOI22_X1 port map( A1 => REGISTERS_24_49_port, A2 => n365, B1 => 
                           REGISTERS_26_49_port, B2 => n328, ZN => n1960);
   U2031 : AND4_X1 port map( A1 => n1963, A2 => n1962, A3 => n1961, A4 => n1960
                           , ZN => n1975);
   U2032 : AOI22_X1 port map( A1 => REGISTERS_5_49_port, A2 => n143_port, B1 =>
                           REGISTERS_7_49_port, B2 => n106_port, ZN => n1967);
   U2033 : AOI22_X1 port map( A1 => REGISTERS_1_49_port, A2 => n217, B1 => 
                           REGISTERS_3_49_port, B2 => n180, ZN => n1966);
   U2034 : AOI22_X1 port map( A1 => REGISTERS_4_49_port, A2 => n291, B1 => 
                           REGISTERS_6_49_port, B2 => n254_port, ZN => n1965);
   U2035 : AOI22_X1 port map( A1 => REGISTERS_0_49_port, A2 => n365, B1 => 
                           REGISTERS_2_49_port, B2 => n328, ZN => n1964);
   U2036 : NAND4_X1 port map( A1 => n1967, A2 => n1966, A3 => n1965, A4 => 
                           n1964, ZN => n1973);
   U2037 : AOI22_X1 port map( A1 => REGISTERS_13_49_port, A2 => n143_port, B1 
                           => REGISTERS_15_49_port, B2 => n106_port, ZN => 
                           n1971);
   U2038 : AOI22_X1 port map( A1 => REGISTERS_9_49_port, A2 => n217, B1 => 
                           REGISTERS_11_49_port, B2 => n180, ZN => n1970);
   U2039 : AOI22_X1 port map( A1 => REGISTERS_12_49_port, A2 => n291, B1 => 
                           REGISTERS_14_49_port, B2 => n254_port, ZN => n1969);
   U2040 : AOI22_X1 port map( A1 => REGISTERS_8_49_port, A2 => n365, B1 => 
                           REGISTERS_10_49_port, B2 => n328, ZN => n1968);
   U2041 : NAND4_X1 port map( A1 => n1971, A2 => n1970, A3 => n1969, A4 => 
                           n1968, ZN => n1972);
   U2042 : AOI22_X1 port map( A1 => n1973, A2 => n27, B1 => n1972, B2 => n24, 
                           ZN => n1974);
   U2043 : OAI221_X1 port map( B1 => n2271, B2 => n1976, C1 => n2269, C2 => 
                           n1975, A => n1974, ZN => N110);
   U2044 : AOI22_X1 port map( A1 => REGISTERS_21_50_port, A2 => n143_port, B1 
                           => REGISTERS_23_50_port, B2 => n106_port, ZN => 
                           n1980);
   U2045 : AOI22_X1 port map( A1 => REGISTERS_17_50_port, A2 => n217, B1 => 
                           REGISTERS_19_50_port, B2 => n180, ZN => n1979);
   U2046 : AOI22_X1 port map( A1 => REGISTERS_20_50_port, A2 => n291, B1 => 
                           REGISTERS_22_50_port, B2 => n254_port, ZN => n1978);
   U2047 : AOI22_X1 port map( A1 => REGISTERS_16_50_port, A2 => n365, B1 => 
                           REGISTERS_18_50_port, B2 => n328, ZN => n1977);
   U2048 : AND4_X1 port map( A1 => n1980, A2 => n1979, A3 => n1978, A4 => n1977
                           , ZN => n1997);
   U2049 : AOI22_X1 port map( A1 => REGISTERS_29_50_port, A2 => n143_port, B1 
                           => REGISTERS_31_50_port, B2 => n106_port, ZN => 
                           n1984);
   U2050 : AOI22_X1 port map( A1 => REGISTERS_25_50_port, A2 => n217, B1 => 
                           REGISTERS_27_50_port, B2 => n180, ZN => n1983);
   U2051 : AOI22_X1 port map( A1 => REGISTERS_28_50_port, A2 => n291, B1 => 
                           REGISTERS_30_50_port, B2 => n254_port, ZN => n1982);
   U2052 : AOI22_X1 port map( A1 => REGISTERS_24_50_port, A2 => n365, B1 => 
                           REGISTERS_26_50_port, B2 => n328, ZN => n1981);
   U2053 : AND4_X1 port map( A1 => n1984, A2 => n1983, A3 => n1982, A4 => n1981
                           , ZN => n1996);
   U2054 : AOI22_X1 port map( A1 => REGISTERS_5_50_port, A2 => n143_port, B1 =>
                           REGISTERS_7_50_port, B2 => n106_port, ZN => n1988);
   U2055 : AOI22_X1 port map( A1 => REGISTERS_1_50_port, A2 => n217, B1 => 
                           REGISTERS_3_50_port, B2 => n180, ZN => n1987);
   U2056 : AOI22_X1 port map( A1 => REGISTERS_4_50_port, A2 => n291, B1 => 
                           REGISTERS_6_50_port, B2 => n254_port, ZN => n1986);
   U2057 : AOI22_X1 port map( A1 => REGISTERS_0_50_port, A2 => n365, B1 => 
                           REGISTERS_2_50_port, B2 => n328, ZN => n1985);
   U2058 : NAND4_X1 port map( A1 => n1988, A2 => n1987, A3 => n1986, A4 => 
                           n1985, ZN => n1994);
   U2059 : AOI22_X1 port map( A1 => REGISTERS_13_50_port, A2 => n143_port, B1 
                           => REGISTERS_15_50_port, B2 => n106_port, ZN => 
                           n1992);
   U2060 : AOI22_X1 port map( A1 => REGISTERS_9_50_port, A2 => n217, B1 => 
                           REGISTERS_11_50_port, B2 => n180, ZN => n1991);
   U2061 : AOI22_X1 port map( A1 => REGISTERS_12_50_port, A2 => n291, B1 => 
                           REGISTERS_14_50_port, B2 => n254_port, ZN => n1990);
   U2062 : AOI22_X1 port map( A1 => REGISTERS_8_50_port, A2 => n365, B1 => 
                           REGISTERS_10_50_port, B2 => n328, ZN => n1989);
   U2063 : NAND4_X1 port map( A1 => n1992, A2 => n1991, A3 => n1990, A4 => 
                           n1989, ZN => n1993);
   U2064 : AOI22_X1 port map( A1 => n1994, A2 => n27, B1 => n1993, B2 => n24, 
                           ZN => n1995);
   U2065 : OAI221_X1 port map( B1 => n2271, B2 => n1997, C1 => n2269, C2 => 
                           n1996, A => n1995, ZN => N109);
   U2066 : AOI22_X1 port map( A1 => REGISTERS_21_51_port, A2 => n144_port, B1 
                           => REGISTERS_23_51_port, B2 => n107_port, ZN => 
                           n2001);
   U2067 : AOI22_X1 port map( A1 => REGISTERS_17_51_port, A2 => n218, B1 => 
                           REGISTERS_19_51_port, B2 => n181, ZN => n2000);
   U2068 : AOI22_X1 port map( A1 => REGISTERS_20_51_port, A2 => n292, B1 => 
                           REGISTERS_22_51_port, B2 => n255_port, ZN => n1999);
   U2069 : AOI22_X1 port map( A1 => REGISTERS_16_51_port, A2 => n366, B1 => 
                           REGISTERS_18_51_port, B2 => n329, ZN => n1998);
   U2070 : AND4_X1 port map( A1 => n2001, A2 => n2000, A3 => n1999, A4 => n1998
                           , ZN => n2018);
   U2071 : AOI22_X1 port map( A1 => REGISTERS_29_51_port, A2 => n144_port, B1 
                           => REGISTERS_31_51_port, B2 => n107_port, ZN => 
                           n2005);
   U2072 : AOI22_X1 port map( A1 => REGISTERS_25_51_port, A2 => n218, B1 => 
                           REGISTERS_27_51_port, B2 => n181, ZN => n2004);
   U2073 : AOI22_X1 port map( A1 => REGISTERS_28_51_port, A2 => n292, B1 => 
                           REGISTERS_30_51_port, B2 => n255_port, ZN => n2003);
   U2074 : AOI22_X1 port map( A1 => REGISTERS_24_51_port, A2 => n366, B1 => 
                           REGISTERS_26_51_port, B2 => n329, ZN => n2002);
   U2075 : AND4_X1 port map( A1 => n2005, A2 => n2004, A3 => n2003, A4 => n2002
                           , ZN => n2017);
   U2076 : AOI22_X1 port map( A1 => REGISTERS_5_51_port, A2 => n144_port, B1 =>
                           REGISTERS_7_51_port, B2 => n107_port, ZN => n2009);
   U2077 : AOI22_X1 port map( A1 => REGISTERS_1_51_port, A2 => n218, B1 => 
                           REGISTERS_3_51_port, B2 => n181, ZN => n2008);
   U2078 : AOI22_X1 port map( A1 => REGISTERS_4_51_port, A2 => n292, B1 => 
                           REGISTERS_6_51_port, B2 => n255_port, ZN => n2007);
   U2079 : AOI22_X1 port map( A1 => REGISTERS_0_51_port, A2 => n366, B1 => 
                           REGISTERS_2_51_port, B2 => n329, ZN => n2006);
   U2080 : NAND4_X1 port map( A1 => n2009, A2 => n2008, A3 => n2007, A4 => 
                           n2006, ZN => n2015);
   U2081 : AOI22_X1 port map( A1 => REGISTERS_13_51_port, A2 => n144_port, B1 
                           => REGISTERS_15_51_port, B2 => n107_port, ZN => 
                           n2013);
   U2082 : AOI22_X1 port map( A1 => REGISTERS_9_51_port, A2 => n218, B1 => 
                           REGISTERS_11_51_port, B2 => n181, ZN => n2012);
   U2083 : AOI22_X1 port map( A1 => REGISTERS_12_51_port, A2 => n292, B1 => 
                           REGISTERS_14_51_port, B2 => n255_port, ZN => n2011);
   U2084 : AOI22_X1 port map( A1 => REGISTERS_8_51_port, A2 => n366, B1 => 
                           REGISTERS_10_51_port, B2 => n329, ZN => n2010);
   U2085 : NAND4_X1 port map( A1 => n2013, A2 => n2012, A3 => n2011, A4 => 
                           n2010, ZN => n2014);
   U2086 : AOI22_X1 port map( A1 => n2015, A2 => n27, B1 => n2014, B2 => n24, 
                           ZN => n2016);
   U2087 : OAI221_X1 port map( B1 => n2271, B2 => n2018, C1 => n2269, C2 => 
                           n2017, A => n2016, ZN => N108);
   U2088 : AOI22_X1 port map( A1 => REGISTERS_21_52_port, A2 => n144_port, B1 
                           => REGISTERS_23_52_port, B2 => n107_port, ZN => 
                           n2022);
   U2089 : AOI22_X1 port map( A1 => REGISTERS_17_52_port, A2 => n218, B1 => 
                           REGISTERS_19_52_port, B2 => n181, ZN => n2021);
   U2090 : AOI22_X1 port map( A1 => REGISTERS_20_52_port, A2 => n292, B1 => 
                           REGISTERS_22_52_port, B2 => n255_port, ZN => n2020);
   U2091 : AOI22_X1 port map( A1 => REGISTERS_16_52_port, A2 => n366, B1 => 
                           REGISTERS_18_52_port, B2 => n329, ZN => n2019);
   U2092 : AND4_X1 port map( A1 => n2022, A2 => n2021, A3 => n2020, A4 => n2019
                           , ZN => n2039);
   U2093 : AOI22_X1 port map( A1 => REGISTERS_29_52_port, A2 => n144_port, B1 
                           => REGISTERS_31_52_port, B2 => n107_port, ZN => 
                           n2026);
   U2094 : AOI22_X1 port map( A1 => REGISTERS_25_52_port, A2 => n218, B1 => 
                           REGISTERS_27_52_port, B2 => n181, ZN => n2025);
   U2095 : AOI22_X1 port map( A1 => REGISTERS_28_52_port, A2 => n292, B1 => 
                           REGISTERS_30_52_port, B2 => n255_port, ZN => n2024);
   U2096 : AOI22_X1 port map( A1 => REGISTERS_24_52_port, A2 => n366, B1 => 
                           REGISTERS_26_52_port, B2 => n329, ZN => n2023);
   U2097 : AND4_X1 port map( A1 => n2026, A2 => n2025, A3 => n2024, A4 => n2023
                           , ZN => n2038);
   U2098 : AOI22_X1 port map( A1 => REGISTERS_5_52_port, A2 => n144_port, B1 =>
                           REGISTERS_7_52_port, B2 => n107_port, ZN => n2030);
   U2099 : AOI22_X1 port map( A1 => REGISTERS_1_52_port, A2 => n218, B1 => 
                           REGISTERS_3_52_port, B2 => n181, ZN => n2029);
   U2100 : AOI22_X1 port map( A1 => REGISTERS_4_52_port, A2 => n292, B1 => 
                           REGISTERS_6_52_port, B2 => n255_port, ZN => n2028);
   U2101 : AOI22_X1 port map( A1 => REGISTERS_0_52_port, A2 => n366, B1 => 
                           REGISTERS_2_52_port, B2 => n329, ZN => n2027);
   U2102 : NAND4_X1 port map( A1 => n2030, A2 => n2029, A3 => n2028, A4 => 
                           n2027, ZN => n2036);
   U2103 : AOI22_X1 port map( A1 => REGISTERS_13_52_port, A2 => n144_port, B1 
                           => REGISTERS_15_52_port, B2 => n107_port, ZN => 
                           n2034);
   U2104 : AOI22_X1 port map( A1 => REGISTERS_9_52_port, A2 => n218, B1 => 
                           REGISTERS_11_52_port, B2 => n181, ZN => n2033);
   U2105 : AOI22_X1 port map( A1 => REGISTERS_12_52_port, A2 => n292, B1 => 
                           REGISTERS_14_52_port, B2 => n255_port, ZN => n2032);
   U2106 : AOI22_X1 port map( A1 => REGISTERS_8_52_port, A2 => n366, B1 => 
                           REGISTERS_10_52_port, B2 => n329, ZN => n2031);
   U2107 : NAND4_X1 port map( A1 => n2034, A2 => n2033, A3 => n2032, A4 => 
                           n2031, ZN => n2035);
   U2108 : AOI22_X1 port map( A1 => n2036, A2 => n27, B1 => n2035, B2 => n24, 
                           ZN => n2037);
   U2109 : OAI221_X1 port map( B1 => n2271, B2 => n2039, C1 => n2269, C2 => 
                           n2038, A => n2037, ZN => N107);
   U2110 : AOI22_X1 port map( A1 => REGISTERS_21_53_port, A2 => n144_port, B1 
                           => REGISTERS_23_53_port, B2 => n107_port, ZN => 
                           n2043);
   U2111 : AOI22_X1 port map( A1 => REGISTERS_17_53_port, A2 => n218, B1 => 
                           REGISTERS_19_53_port, B2 => n181, ZN => n2042);
   U2112 : AOI22_X1 port map( A1 => REGISTERS_20_53_port, A2 => n292, B1 => 
                           REGISTERS_22_53_port, B2 => n255_port, ZN => n2041);
   U2113 : AOI22_X1 port map( A1 => REGISTERS_16_53_port, A2 => n366, B1 => 
                           REGISTERS_18_53_port, B2 => n329, ZN => n2040);
   U2114 : AND4_X1 port map( A1 => n2043, A2 => n2042, A3 => n2041, A4 => n2040
                           , ZN => n2060);
   U2115 : AOI22_X1 port map( A1 => REGISTERS_29_53_port, A2 => n144_port, B1 
                           => REGISTERS_31_53_port, B2 => n107_port, ZN => 
                           n2047);
   U2116 : AOI22_X1 port map( A1 => REGISTERS_25_53_port, A2 => n218, B1 => 
                           REGISTERS_27_53_port, B2 => n181, ZN => n2046);
   U2117 : AOI22_X1 port map( A1 => REGISTERS_28_53_port, A2 => n292, B1 => 
                           REGISTERS_30_53_port, B2 => n255_port, ZN => n2045);
   U2118 : AOI22_X1 port map( A1 => REGISTERS_24_53_port, A2 => n366, B1 => 
                           REGISTERS_26_53_port, B2 => n329, ZN => n2044);
   U2119 : AND4_X1 port map( A1 => n2047, A2 => n2046, A3 => n2045, A4 => n2044
                           , ZN => n2059);
   U2120 : AOI22_X1 port map( A1 => REGISTERS_5_53_port, A2 => n144_port, B1 =>
                           REGISTERS_7_53_port, B2 => n107_port, ZN => n2051);
   U2121 : AOI22_X1 port map( A1 => REGISTERS_1_53_port, A2 => n218, B1 => 
                           REGISTERS_3_53_port, B2 => n181, ZN => n2050);
   U2122 : AOI22_X1 port map( A1 => REGISTERS_4_53_port, A2 => n292, B1 => 
                           REGISTERS_6_53_port, B2 => n255_port, ZN => n2049);
   U2123 : AOI22_X1 port map( A1 => REGISTERS_0_53_port, A2 => n366, B1 => 
                           REGISTERS_2_53_port, B2 => n329, ZN => n2048);
   U2124 : NAND4_X1 port map( A1 => n2051, A2 => n2050, A3 => n2049, A4 => 
                           n2048, ZN => n2057);
   U2125 : AOI22_X1 port map( A1 => REGISTERS_13_53_port, A2 => n144_port, B1 
                           => REGISTERS_15_53_port, B2 => n107_port, ZN => 
                           n2055);
   U2126 : AOI22_X1 port map( A1 => REGISTERS_9_53_port, A2 => n218, B1 => 
                           REGISTERS_11_53_port, B2 => n181, ZN => n2054);
   U2127 : AOI22_X1 port map( A1 => REGISTERS_12_53_port, A2 => n292, B1 => 
                           REGISTERS_14_53_port, B2 => n255_port, ZN => n2053);
   U2128 : AOI22_X1 port map( A1 => REGISTERS_8_53_port, A2 => n366, B1 => 
                           REGISTERS_10_53_port, B2 => n329, ZN => n2052);
   U2129 : NAND4_X1 port map( A1 => n2055, A2 => n2054, A3 => n2053, A4 => 
                           n2052, ZN => n2056);
   U2130 : AOI22_X1 port map( A1 => n2057, A2 => n27, B1 => n2056, B2 => n24, 
                           ZN => n2058);
   U2131 : OAI221_X1 port map( B1 => n2271, B2 => n2060, C1 => n2269, C2 => 
                           n2059, A => n2058, ZN => N106);
   U2132 : AOI22_X1 port map( A1 => REGISTERS_21_54_port, A2 => n145_port, B1 
                           => REGISTERS_23_54_port, B2 => n108_port, ZN => 
                           n2064);
   U2133 : AOI22_X1 port map( A1 => REGISTERS_17_54_port, A2 => n219, B1 => 
                           REGISTERS_19_54_port, B2 => n182, ZN => n2063);
   U2134 : AOI22_X1 port map( A1 => REGISTERS_20_54_port, A2 => n293, B1 => 
                           REGISTERS_22_54_port, B2 => n256_port, ZN => n2062);
   U2135 : AOI22_X1 port map( A1 => REGISTERS_16_54_port, A2 => n367, B1 => 
                           REGISTERS_18_54_port, B2 => n330, ZN => n2061);
   U2136 : AND4_X1 port map( A1 => n2064, A2 => n2063, A3 => n2062, A4 => n2061
                           , ZN => n2081);
   U2137 : AOI22_X1 port map( A1 => REGISTERS_29_54_port, A2 => n145_port, B1 
                           => REGISTERS_31_54_port, B2 => n108_port, ZN => 
                           n2068);
   U2138 : AOI22_X1 port map( A1 => REGISTERS_25_54_port, A2 => n219, B1 => 
                           REGISTERS_27_54_port, B2 => n182, ZN => n2067);
   U2139 : AOI22_X1 port map( A1 => REGISTERS_28_54_port, A2 => n293, B1 => 
                           REGISTERS_30_54_port, B2 => n256_port, ZN => n2066);
   U2140 : AOI22_X1 port map( A1 => REGISTERS_24_54_port, A2 => n367, B1 => 
                           REGISTERS_26_54_port, B2 => n330, ZN => n2065);
   U2141 : AND4_X1 port map( A1 => n2068, A2 => n2067, A3 => n2066, A4 => n2065
                           , ZN => n2080);
   U2142 : AOI22_X1 port map( A1 => REGISTERS_5_54_port, A2 => n145_port, B1 =>
                           REGISTERS_7_54_port, B2 => n108_port, ZN => n2072);
   U2143 : AOI22_X1 port map( A1 => REGISTERS_1_54_port, A2 => n219, B1 => 
                           REGISTERS_3_54_port, B2 => n182, ZN => n2071);
   U2144 : AOI22_X1 port map( A1 => REGISTERS_4_54_port, A2 => n293, B1 => 
                           REGISTERS_6_54_port, B2 => n256_port, ZN => n2070);
   U2145 : AOI22_X1 port map( A1 => REGISTERS_0_54_port, A2 => n367, B1 => 
                           REGISTERS_2_54_port, B2 => n330, ZN => n2069);
   U2146 : NAND4_X1 port map( A1 => n2072, A2 => n2071, A3 => n2070, A4 => 
                           n2069, ZN => n2078);
   U2147 : AOI22_X1 port map( A1 => REGISTERS_13_54_port, A2 => n145_port, B1 
                           => REGISTERS_15_54_port, B2 => n108_port, ZN => 
                           n2076);
   U2148 : AOI22_X1 port map( A1 => REGISTERS_9_54_port, A2 => n219, B1 => 
                           REGISTERS_11_54_port, B2 => n182, ZN => n2075);
   U2149 : AOI22_X1 port map( A1 => REGISTERS_12_54_port, A2 => n293, B1 => 
                           REGISTERS_14_54_port, B2 => n256_port, ZN => n2074);
   U2150 : AOI22_X1 port map( A1 => REGISTERS_8_54_port, A2 => n367, B1 => 
                           REGISTERS_10_54_port, B2 => n330, ZN => n2073);
   U2151 : NAND4_X1 port map( A1 => n2076, A2 => n2075, A3 => n2074, A4 => 
                           n2073, ZN => n2077);
   U2152 : AOI22_X1 port map( A1 => n2078, A2 => n27, B1 => n2077, B2 => n24, 
                           ZN => n2079);
   U2153 : OAI221_X1 port map( B1 => n2271, B2 => n2081, C1 => n2269, C2 => 
                           n2080, A => n2079, ZN => N105);
   U2154 : AOI22_X1 port map( A1 => REGISTERS_21_55_port, A2 => n145_port, B1 
                           => REGISTERS_23_55_port, B2 => n108_port, ZN => 
                           n2085);
   U2155 : AOI22_X1 port map( A1 => REGISTERS_17_55_port, A2 => n219, B1 => 
                           REGISTERS_19_55_port, B2 => n182, ZN => n2084);
   U2156 : AOI22_X1 port map( A1 => REGISTERS_20_55_port, A2 => n293, B1 => 
                           REGISTERS_22_55_port, B2 => n256_port, ZN => n2083);
   U2157 : AOI22_X1 port map( A1 => REGISTERS_16_55_port, A2 => n367, B1 => 
                           REGISTERS_18_55_port, B2 => n330, ZN => n2082);
   U2158 : AND4_X1 port map( A1 => n2085, A2 => n2084, A3 => n2083, A4 => n2082
                           , ZN => n2102);
   U2159 : AOI22_X1 port map( A1 => REGISTERS_29_55_port, A2 => n145_port, B1 
                           => REGISTERS_31_55_port, B2 => n108_port, ZN => 
                           n2089);
   U2160 : AOI22_X1 port map( A1 => REGISTERS_25_55_port, A2 => n219, B1 => 
                           REGISTERS_27_55_port, B2 => n182, ZN => n2088);
   U2161 : AOI22_X1 port map( A1 => REGISTERS_28_55_port, A2 => n293, B1 => 
                           REGISTERS_30_55_port, B2 => n256_port, ZN => n2087);
   U2162 : AOI22_X1 port map( A1 => REGISTERS_24_55_port, A2 => n367, B1 => 
                           REGISTERS_26_55_port, B2 => n330, ZN => n2086);
   U2163 : AND4_X1 port map( A1 => n2089, A2 => n2088, A3 => n2087, A4 => n2086
                           , ZN => n2101);
   U2164 : AOI22_X1 port map( A1 => REGISTERS_5_55_port, A2 => n145_port, B1 =>
                           REGISTERS_7_55_port, B2 => n108_port, ZN => n2093);
   U2165 : AOI22_X1 port map( A1 => REGISTERS_1_55_port, A2 => n219, B1 => 
                           REGISTERS_3_55_port, B2 => n182, ZN => n2092);
   U2166 : AOI22_X1 port map( A1 => REGISTERS_4_55_port, A2 => n293, B1 => 
                           REGISTERS_6_55_port, B2 => n256_port, ZN => n2091);
   U2167 : AOI22_X1 port map( A1 => REGISTERS_0_55_port, A2 => n367, B1 => 
                           REGISTERS_2_55_port, B2 => n330, ZN => n2090);
   U2168 : NAND4_X1 port map( A1 => n2093, A2 => n2092, A3 => n2091, A4 => 
                           n2090, ZN => n2099);
   U2169 : AOI22_X1 port map( A1 => REGISTERS_13_55_port, A2 => n145_port, B1 
                           => REGISTERS_15_55_port, B2 => n108_port, ZN => 
                           n2097);
   U2170 : AOI22_X1 port map( A1 => REGISTERS_9_55_port, A2 => n219, B1 => 
                           REGISTERS_11_55_port, B2 => n182, ZN => n2096);
   U2171 : AOI22_X1 port map( A1 => REGISTERS_12_55_port, A2 => n293, B1 => 
                           REGISTERS_14_55_port, B2 => n256_port, ZN => n2095);
   U2172 : AOI22_X1 port map( A1 => REGISTERS_8_55_port, A2 => n367, B1 => 
                           REGISTERS_10_55_port, B2 => n330, ZN => n2094);
   U2173 : NAND4_X1 port map( A1 => n2097, A2 => n2096, A3 => n2095, A4 => 
                           n2094, ZN => n2098);
   U2174 : AOI22_X1 port map( A1 => n2099, A2 => n27, B1 => n2098, B2 => n24, 
                           ZN => n2100);
   U2175 : OAI221_X1 port map( B1 => n2271, B2 => n2102, C1 => n2269, C2 => 
                           n2101, A => n2100, ZN => N104);
   U2176 : AOI22_X1 port map( A1 => REGISTERS_21_56_port, A2 => n145_port, B1 
                           => REGISTERS_23_56_port, B2 => n108_port, ZN => 
                           n2106);
   U2177 : AOI22_X1 port map( A1 => REGISTERS_17_56_port, A2 => n219, B1 => 
                           REGISTERS_19_56_port, B2 => n182, ZN => n2105);
   U2178 : AOI22_X1 port map( A1 => REGISTERS_20_56_port, A2 => n293, B1 => 
                           REGISTERS_22_56_port, B2 => n256_port, ZN => n2104);
   U2179 : AOI22_X1 port map( A1 => REGISTERS_16_56_port, A2 => n367, B1 => 
                           REGISTERS_18_56_port, B2 => n330, ZN => n2103);
   U2180 : AND4_X1 port map( A1 => n2106, A2 => n2105, A3 => n2104, A4 => n2103
                           , ZN => n2123);
   U2181 : AOI22_X1 port map( A1 => REGISTERS_29_56_port, A2 => n145_port, B1 
                           => REGISTERS_31_56_port, B2 => n108_port, ZN => 
                           n2110);
   U2182 : AOI22_X1 port map( A1 => REGISTERS_25_56_port, A2 => n219, B1 => 
                           REGISTERS_27_56_port, B2 => n182, ZN => n2109);
   U2183 : AOI22_X1 port map( A1 => REGISTERS_28_56_port, A2 => n293, B1 => 
                           REGISTERS_30_56_port, B2 => n256_port, ZN => n2108);
   U2184 : AOI22_X1 port map( A1 => REGISTERS_24_56_port, A2 => n367, B1 => 
                           REGISTERS_26_56_port, B2 => n330, ZN => n2107);
   U2185 : AND4_X1 port map( A1 => n2110, A2 => n2109, A3 => n2108, A4 => n2107
                           , ZN => n2122);
   U2186 : AOI22_X1 port map( A1 => REGISTERS_5_56_port, A2 => n145_port, B1 =>
                           REGISTERS_7_56_port, B2 => n108_port, ZN => n2114);
   U2187 : AOI22_X1 port map( A1 => REGISTERS_1_56_port, A2 => n219, B1 => 
                           REGISTERS_3_56_port, B2 => n182, ZN => n2113);
   U2188 : AOI22_X1 port map( A1 => REGISTERS_4_56_port, A2 => n293, B1 => 
                           REGISTERS_6_56_port, B2 => n256_port, ZN => n2112);
   U2189 : AOI22_X1 port map( A1 => REGISTERS_0_56_port, A2 => n367, B1 => 
                           REGISTERS_2_56_port, B2 => n330, ZN => n2111);
   U2190 : NAND4_X1 port map( A1 => n2114, A2 => n2113, A3 => n2112, A4 => 
                           n2111, ZN => n2120);
   U2191 : AOI22_X1 port map( A1 => REGISTERS_13_56_port, A2 => n145_port, B1 
                           => REGISTERS_15_56_port, B2 => n108_port, ZN => 
                           n2118);
   U2192 : AOI22_X1 port map( A1 => REGISTERS_9_56_port, A2 => n219, B1 => 
                           REGISTERS_11_56_port, B2 => n182, ZN => n2117);
   U2193 : AOI22_X1 port map( A1 => REGISTERS_12_56_port, A2 => n293, B1 => 
                           REGISTERS_14_56_port, B2 => n256_port, ZN => n2116);
   U2194 : AOI22_X1 port map( A1 => REGISTERS_8_56_port, A2 => n367, B1 => 
                           REGISTERS_10_56_port, B2 => n330, ZN => n2115);
   U2195 : NAND4_X1 port map( A1 => n2118, A2 => n2117, A3 => n2116, A4 => 
                           n2115, ZN => n2119);
   U2196 : AOI22_X1 port map( A1 => n2120, A2 => n27, B1 => n2119, B2 => n24, 
                           ZN => n2121);
   U2197 : OAI221_X1 port map( B1 => n2271, B2 => n2123, C1 => n2269, C2 => 
                           n2122, A => n2121, ZN => N103);
   U2198 : AOI22_X1 port map( A1 => REGISTERS_21_57_port, A2 => n146_port, B1 
                           => REGISTERS_23_57_port, B2 => n109_port, ZN => 
                           n2127);
   U2199 : AOI22_X1 port map( A1 => REGISTERS_17_57_port, A2 => n220, B1 => 
                           REGISTERS_19_57_port, B2 => n183, ZN => n2126);
   U2200 : AOI22_X1 port map( A1 => REGISTERS_20_57_port, A2 => n294, B1 => 
                           REGISTERS_22_57_port, B2 => n257_port, ZN => n2125);
   U2201 : AOI22_X1 port map( A1 => REGISTERS_16_57_port, A2 => n368, B1 => 
                           REGISTERS_18_57_port, B2 => n331, ZN => n2124);
   U2202 : AND4_X1 port map( A1 => n2127, A2 => n2126, A3 => n2125, A4 => n2124
                           , ZN => n2144);
   U2203 : AOI22_X1 port map( A1 => REGISTERS_29_57_port, A2 => n146_port, B1 
                           => REGISTERS_31_57_port, B2 => n109_port, ZN => 
                           n2131);
   U2204 : AOI22_X1 port map( A1 => REGISTERS_25_57_port, A2 => n220, B1 => 
                           REGISTERS_27_57_port, B2 => n183, ZN => n2130);
   U2205 : AOI22_X1 port map( A1 => REGISTERS_28_57_port, A2 => n294, B1 => 
                           REGISTERS_30_57_port, B2 => n257_port, ZN => n2129);
   U2206 : AOI22_X1 port map( A1 => REGISTERS_24_57_port, A2 => n368, B1 => 
                           REGISTERS_26_57_port, B2 => n331, ZN => n2128);
   U2207 : AND4_X1 port map( A1 => n2131, A2 => n2130, A3 => n2129, A4 => n2128
                           , ZN => n2143);
   U2208 : AOI22_X1 port map( A1 => REGISTERS_5_57_port, A2 => n146_port, B1 =>
                           REGISTERS_7_57_port, B2 => n109_port, ZN => n2135);
   U2209 : AOI22_X1 port map( A1 => REGISTERS_1_57_port, A2 => n220, B1 => 
                           REGISTERS_3_57_port, B2 => n183, ZN => n2134);
   U2210 : AOI22_X1 port map( A1 => REGISTERS_4_57_port, A2 => n294, B1 => 
                           REGISTERS_6_57_port, B2 => n257_port, ZN => n2133);
   U2211 : AOI22_X1 port map( A1 => REGISTERS_0_57_port, A2 => n368, B1 => 
                           REGISTERS_2_57_port, B2 => n331, ZN => n2132);
   U2212 : NAND4_X1 port map( A1 => n2135, A2 => n2134, A3 => n2133, A4 => 
                           n2132, ZN => n2141);
   U2213 : AOI22_X1 port map( A1 => REGISTERS_13_57_port, A2 => n146_port, B1 
                           => REGISTERS_15_57_port, B2 => n109_port, ZN => 
                           n2139);
   U2214 : AOI22_X1 port map( A1 => REGISTERS_9_57_port, A2 => n220, B1 => 
                           REGISTERS_11_57_port, B2 => n183, ZN => n2138);
   U2215 : AOI22_X1 port map( A1 => REGISTERS_12_57_port, A2 => n294, B1 => 
                           REGISTERS_14_57_port, B2 => n257_port, ZN => n2137);
   U2216 : AOI22_X1 port map( A1 => REGISTERS_8_57_port, A2 => n368, B1 => 
                           REGISTERS_10_57_port, B2 => n331, ZN => n2136);
   U2217 : NAND4_X1 port map( A1 => n2139, A2 => n2138, A3 => n2137, A4 => 
                           n2136, ZN => n2140);
   U2218 : AOI22_X1 port map( A1 => n2141, A2 => n27, B1 => n2140, B2 => n24, 
                           ZN => n2142);
   U2219 : OAI221_X1 port map( B1 => n2271, B2 => n2144, C1 => n2269, C2 => 
                           n2143, A => n2142, ZN => N102);
   U2220 : AOI22_X1 port map( A1 => REGISTERS_21_58_port, A2 => n146_port, B1 
                           => REGISTERS_23_58_port, B2 => n109_port, ZN => 
                           n2148);
   U2221 : AOI22_X1 port map( A1 => REGISTERS_17_58_port, A2 => n220, B1 => 
                           REGISTERS_19_58_port, B2 => n183, ZN => n2147);
   U2222 : AOI22_X1 port map( A1 => REGISTERS_20_58_port, A2 => n294, B1 => 
                           REGISTERS_22_58_port, B2 => n257_port, ZN => n2146);
   U2223 : AOI22_X1 port map( A1 => REGISTERS_16_58_port, A2 => n368, B1 => 
                           REGISTERS_18_58_port, B2 => n331, ZN => n2145);
   U2224 : AND4_X1 port map( A1 => n2148, A2 => n2147, A3 => n2146, A4 => n2145
                           , ZN => n2165);
   U2225 : AOI22_X1 port map( A1 => REGISTERS_29_58_port, A2 => n146_port, B1 
                           => REGISTERS_31_58_port, B2 => n109_port, ZN => 
                           n2152);
   U2226 : AOI22_X1 port map( A1 => REGISTERS_25_58_port, A2 => n220, B1 => 
                           REGISTERS_27_58_port, B2 => n183, ZN => n2151);
   U2227 : AOI22_X1 port map( A1 => REGISTERS_28_58_port, A2 => n294, B1 => 
                           REGISTERS_30_58_port, B2 => n257_port, ZN => n2150);
   U2228 : AOI22_X1 port map( A1 => REGISTERS_24_58_port, A2 => n368, B1 => 
                           REGISTERS_26_58_port, B2 => n331, ZN => n2149);
   U2229 : AND4_X1 port map( A1 => n2152, A2 => n2151, A3 => n2150, A4 => n2149
                           , ZN => n2164);
   U2230 : AOI22_X1 port map( A1 => REGISTERS_5_58_port, A2 => n146_port, B1 =>
                           REGISTERS_7_58_port, B2 => n109_port, ZN => n2156);
   U2231 : AOI22_X1 port map( A1 => REGISTERS_1_58_port, A2 => n220, B1 => 
                           REGISTERS_3_58_port, B2 => n183, ZN => n2155);
   U2232 : AOI22_X1 port map( A1 => REGISTERS_4_58_port, A2 => n294, B1 => 
                           REGISTERS_6_58_port, B2 => n257_port, ZN => n2154);
   U2233 : AOI22_X1 port map( A1 => REGISTERS_0_58_port, A2 => n368, B1 => 
                           REGISTERS_2_58_port, B2 => n331, ZN => n2153);
   U2234 : NAND4_X1 port map( A1 => n2156, A2 => n2155, A3 => n2154, A4 => 
                           n2153, ZN => n2162);
   U2235 : AOI22_X1 port map( A1 => REGISTERS_13_58_port, A2 => n146_port, B1 
                           => REGISTERS_15_58_port, B2 => n109_port, ZN => 
                           n2160);
   U2236 : AOI22_X1 port map( A1 => REGISTERS_9_58_port, A2 => n220, B1 => 
                           REGISTERS_11_58_port, B2 => n183, ZN => n2159);
   U2237 : AOI22_X1 port map( A1 => REGISTERS_12_58_port, A2 => n294, B1 => 
                           REGISTERS_14_58_port, B2 => n257_port, ZN => n2158);
   U2238 : AOI22_X1 port map( A1 => REGISTERS_8_58_port, A2 => n368, B1 => 
                           REGISTERS_10_58_port, B2 => n331, ZN => n2157);
   U2239 : NAND4_X1 port map( A1 => n2160, A2 => n2159, A3 => n2158, A4 => 
                           n2157, ZN => n2161);
   U2240 : AOI22_X1 port map( A1 => n2162, A2 => n27, B1 => n2161, B2 => n24, 
                           ZN => n2163);
   U2241 : OAI221_X1 port map( B1 => n2271, B2 => n2165, C1 => n2269, C2 => 
                           n2164, A => n2163, ZN => N101);
   U2242 : AOI22_X1 port map( A1 => REGISTERS_21_59_port, A2 => n146_port, B1 
                           => REGISTERS_23_59_port, B2 => n109_port, ZN => 
                           n2169);
   U2243 : AOI22_X1 port map( A1 => REGISTERS_17_59_port, A2 => n220, B1 => 
                           REGISTERS_19_59_port, B2 => n183, ZN => n2168);
   U2244 : AOI22_X1 port map( A1 => REGISTERS_20_59_port, A2 => n294, B1 => 
                           REGISTERS_22_59_port, B2 => n257_port, ZN => n2167);
   U2245 : AOI22_X1 port map( A1 => REGISTERS_16_59_port, A2 => n368, B1 => 
                           REGISTERS_18_59_port, B2 => n331, ZN => n2166);
   U2246 : AND4_X1 port map( A1 => n2169, A2 => n2168, A3 => n2167, A4 => n2166
                           , ZN => n2186);
   U2247 : AOI22_X1 port map( A1 => REGISTERS_29_59_port, A2 => n146_port, B1 
                           => REGISTERS_31_59_port, B2 => n109_port, ZN => 
                           n2173);
   U2248 : AOI22_X1 port map( A1 => REGISTERS_25_59_port, A2 => n220, B1 => 
                           REGISTERS_27_59_port, B2 => n183, ZN => n2172);
   U2249 : AOI22_X1 port map( A1 => REGISTERS_28_59_port, A2 => n294, B1 => 
                           REGISTERS_30_59_port, B2 => n257_port, ZN => n2171);
   U2250 : AOI22_X1 port map( A1 => REGISTERS_24_59_port, A2 => n368, B1 => 
                           REGISTERS_26_59_port, B2 => n331, ZN => n2170);
   U2251 : AND4_X1 port map( A1 => n2173, A2 => n2172, A3 => n2171, A4 => n2170
                           , ZN => n2185);
   U2252 : AOI22_X1 port map( A1 => REGISTERS_5_59_port, A2 => n146_port, B1 =>
                           REGISTERS_7_59_port, B2 => n109_port, ZN => n2177);
   U2253 : AOI22_X1 port map( A1 => REGISTERS_1_59_port, A2 => n220, B1 => 
                           REGISTERS_3_59_port, B2 => n183, ZN => n2176);
   U2254 : AOI22_X1 port map( A1 => REGISTERS_4_59_port, A2 => n294, B1 => 
                           REGISTERS_6_59_port, B2 => n257_port, ZN => n2175);
   U2255 : AOI22_X1 port map( A1 => REGISTERS_0_59_port, A2 => n368, B1 => 
                           REGISTERS_2_59_port, B2 => n331, ZN => n2174);
   U2256 : NAND4_X1 port map( A1 => n2177, A2 => n2176, A3 => n2175, A4 => 
                           n2174, ZN => n2183);
   U2257 : AOI22_X1 port map( A1 => REGISTERS_13_59_port, A2 => n146_port, B1 
                           => REGISTERS_15_59_port, B2 => n109_port, ZN => 
                           n2181);
   U2258 : AOI22_X1 port map( A1 => REGISTERS_9_59_port, A2 => n220, B1 => 
                           REGISTERS_11_59_port, B2 => n183, ZN => n2180);
   U2259 : AOI22_X1 port map( A1 => REGISTERS_12_59_port, A2 => n294, B1 => 
                           REGISTERS_14_59_port, B2 => n257_port, ZN => n2179);
   U2260 : AOI22_X1 port map( A1 => REGISTERS_8_59_port, A2 => n368, B1 => 
                           REGISTERS_10_59_port, B2 => n331, ZN => n2178);
   U2261 : NAND4_X1 port map( A1 => n2181, A2 => n2180, A3 => n2179, A4 => 
                           n2178, ZN => n2182);
   U2262 : AOI22_X1 port map( A1 => n2183, A2 => n27, B1 => n2182, B2 => n24, 
                           ZN => n2184);
   U2263 : OAI221_X1 port map( B1 => n2271, B2 => n2186, C1 => n2269, C2 => 
                           n2185, A => n2184, ZN => N100);
   U2264 : AOI22_X1 port map( A1 => REGISTERS_21_60_port, A2 => n147_port, B1 
                           => REGISTERS_23_60_port, B2 => n110_port, ZN => 
                           n2190);
   U2265 : AOI22_X1 port map( A1 => REGISTERS_17_60_port, A2 => n221, B1 => 
                           REGISTERS_19_60_port, B2 => n184, ZN => n2189);
   U2266 : AOI22_X1 port map( A1 => REGISTERS_20_60_port, A2 => n295, B1 => 
                           REGISTERS_22_60_port, B2 => n258_port, ZN => n2188);
   U2267 : AOI22_X1 port map( A1 => REGISTERS_16_60_port, A2 => n369, B1 => 
                           REGISTERS_18_60_port, B2 => n332, ZN => n2187);
   U2268 : AND4_X1 port map( A1 => n2190, A2 => n2189, A3 => n2188, A4 => n2187
                           , ZN => n2207);
   U2269 : AOI22_X1 port map( A1 => REGISTERS_29_60_port, A2 => n147_port, B1 
                           => REGISTERS_31_60_port, B2 => n110_port, ZN => 
                           n2194);
   U2270 : AOI22_X1 port map( A1 => REGISTERS_25_60_port, A2 => n221, B1 => 
                           REGISTERS_27_60_port, B2 => n184, ZN => n2193);
   U2271 : AOI22_X1 port map( A1 => REGISTERS_28_60_port, A2 => n295, B1 => 
                           REGISTERS_30_60_port, B2 => n258_port, ZN => n2192);
   U2272 : AOI22_X1 port map( A1 => REGISTERS_24_60_port, A2 => n369, B1 => 
                           REGISTERS_26_60_port, B2 => n332, ZN => n2191);
   U2273 : AND4_X1 port map( A1 => n2194, A2 => n2193, A3 => n2192, A4 => n2191
                           , ZN => n2206);
   U2274 : AOI22_X1 port map( A1 => REGISTERS_5_60_port, A2 => n147_port, B1 =>
                           REGISTERS_7_60_port, B2 => n110_port, ZN => n2198);
   U2275 : AOI22_X1 port map( A1 => REGISTERS_1_60_port, A2 => n221, B1 => 
                           REGISTERS_3_60_port, B2 => n184, ZN => n2197);
   U2276 : AOI22_X1 port map( A1 => REGISTERS_4_60_port, A2 => n295, B1 => 
                           REGISTERS_6_60_port, B2 => n258_port, ZN => n2196);
   U2277 : AOI22_X1 port map( A1 => REGISTERS_0_60_port, A2 => n369, B1 => 
                           REGISTERS_2_60_port, B2 => n332, ZN => n2195);
   U2278 : NAND4_X1 port map( A1 => n2198, A2 => n2197, A3 => n2196, A4 => 
                           n2195, ZN => n2204);
   U2279 : AOI22_X1 port map( A1 => REGISTERS_13_60_port, A2 => n147_port, B1 
                           => REGISTERS_15_60_port, B2 => n110_port, ZN => 
                           n2202);
   U2280 : AOI22_X1 port map( A1 => REGISTERS_9_60_port, A2 => n221, B1 => 
                           REGISTERS_11_60_port, B2 => n184, ZN => n2201);
   U2281 : AOI22_X1 port map( A1 => REGISTERS_12_60_port, A2 => n295, B1 => 
                           REGISTERS_14_60_port, B2 => n258_port, ZN => n2200);
   U2282 : AOI22_X1 port map( A1 => REGISTERS_8_60_port, A2 => n369, B1 => 
                           REGISTERS_10_60_port, B2 => n332, ZN => n2199);
   U2283 : NAND4_X1 port map( A1 => n2202, A2 => n2201, A3 => n2200, A4 => 
                           n2199, ZN => n2203);
   U2284 : AOI22_X1 port map( A1 => n2204, A2 => n27, B1 => n2203, B2 => n24, 
                           ZN => n2205);
   U2285 : OAI221_X1 port map( B1 => n2271, B2 => n2207, C1 => n2269, C2 => 
                           n2206, A => n2205, ZN => N99);
   U2286 : AOI22_X1 port map( A1 => REGISTERS_21_61_port, A2 => n147_port, B1 
                           => REGISTERS_23_61_port, B2 => n110_port, ZN => 
                           n2211);
   U2287 : AOI22_X1 port map( A1 => REGISTERS_17_61_port, A2 => n221, B1 => 
                           REGISTERS_19_61_port, B2 => n184, ZN => n2210);
   U2288 : AOI22_X1 port map( A1 => REGISTERS_20_61_port, A2 => n295, B1 => 
                           REGISTERS_22_61_port, B2 => n258_port, ZN => n2209);
   U2289 : AOI22_X1 port map( A1 => REGISTERS_16_61_port, A2 => n369, B1 => 
                           REGISTERS_18_61_port, B2 => n332, ZN => n2208);
   U2290 : AND4_X1 port map( A1 => n2211, A2 => n2210, A3 => n2209, A4 => n2208
                           , ZN => n2228);
   U2291 : AOI22_X1 port map( A1 => REGISTERS_29_61_port, A2 => n147_port, B1 
                           => REGISTERS_31_61_port, B2 => n110_port, ZN => 
                           n2215);
   U2292 : AOI22_X1 port map( A1 => REGISTERS_25_61_port, A2 => n221, B1 => 
                           REGISTERS_27_61_port, B2 => n184, ZN => n2214);
   U2293 : AOI22_X1 port map( A1 => REGISTERS_28_61_port, A2 => n295, B1 => 
                           REGISTERS_30_61_port, B2 => n258_port, ZN => n2213);
   U2294 : AOI22_X1 port map( A1 => REGISTERS_24_61_port, A2 => n369, B1 => 
                           REGISTERS_26_61_port, B2 => n332, ZN => n2212);
   U2295 : AND4_X1 port map( A1 => n2215, A2 => n2214, A3 => n2213, A4 => n2212
                           , ZN => n2227);
   U2296 : AOI22_X1 port map( A1 => REGISTERS_5_61_port, A2 => n147_port, B1 =>
                           REGISTERS_7_61_port, B2 => n110_port, ZN => n2219);
   U2297 : AOI22_X1 port map( A1 => REGISTERS_1_61_port, A2 => n221, B1 => 
                           REGISTERS_3_61_port, B2 => n184, ZN => n2218);
   U2298 : AOI22_X1 port map( A1 => REGISTERS_4_61_port, A2 => n295, B1 => 
                           REGISTERS_6_61_port, B2 => n258_port, ZN => n2217);
   U2299 : AOI22_X1 port map( A1 => REGISTERS_0_61_port, A2 => n369, B1 => 
                           REGISTERS_2_61_port, B2 => n332, ZN => n2216);
   U2300 : NAND4_X1 port map( A1 => n2219, A2 => n2218, A3 => n2217, A4 => 
                           n2216, ZN => n2225);
   U2301 : AOI22_X1 port map( A1 => REGISTERS_13_61_port, A2 => n147_port, B1 
                           => REGISTERS_15_61_port, B2 => n110_port, ZN => 
                           n2223);
   U2302 : AOI22_X1 port map( A1 => REGISTERS_9_61_port, A2 => n221, B1 => 
                           REGISTERS_11_61_port, B2 => n184, ZN => n2222);
   U2303 : AOI22_X1 port map( A1 => REGISTERS_12_61_port, A2 => n295, B1 => 
                           REGISTERS_14_61_port, B2 => n258_port, ZN => n2221);
   U2304 : AOI22_X1 port map( A1 => REGISTERS_8_61_port, A2 => n369, B1 => 
                           REGISTERS_10_61_port, B2 => n332, ZN => n2220);
   U2305 : NAND4_X1 port map( A1 => n2223, A2 => n2222, A3 => n2221, A4 => 
                           n2220, ZN => n2224);
   U2306 : AOI22_X1 port map( A1 => n2225, A2 => n27, B1 => n2224, B2 => n24, 
                           ZN => n2226);
   U2307 : OAI221_X1 port map( B1 => n2271, B2 => n2228, C1 => n2269, C2 => 
                           n2227, A => n2226, ZN => N98);
   U2308 : AOI22_X1 port map( A1 => REGISTERS_21_62_port, A2 => n147_port, B1 
                           => REGISTERS_23_62_port, B2 => n110_port, ZN => 
                           n2232);
   U2309 : AOI22_X1 port map( A1 => REGISTERS_17_62_port, A2 => n221, B1 => 
                           REGISTERS_19_62_port, B2 => n184, ZN => n2231);
   U2310 : AOI22_X1 port map( A1 => REGISTERS_20_62_port, A2 => n295, B1 => 
                           REGISTERS_22_62_port, B2 => n258_port, ZN => n2230);
   U2311 : AOI22_X1 port map( A1 => REGISTERS_16_62_port, A2 => n369, B1 => 
                           REGISTERS_18_62_port, B2 => n332, ZN => n2229);
   U2312 : AND4_X1 port map( A1 => n2232, A2 => n2231, A3 => n2230, A4 => n2229
                           , ZN => n2249);
   U2313 : AOI22_X1 port map( A1 => REGISTERS_29_62_port, A2 => n147_port, B1 
                           => REGISTERS_31_62_port, B2 => n110_port, ZN => 
                           n2236);
   U2314 : AOI22_X1 port map( A1 => REGISTERS_25_62_port, A2 => n221, B1 => 
                           REGISTERS_27_62_port, B2 => n184, ZN => n2235);
   U2315 : AOI22_X1 port map( A1 => REGISTERS_28_62_port, A2 => n295, B1 => 
                           REGISTERS_30_62_port, B2 => n258_port, ZN => n2234);
   U2316 : AOI22_X1 port map( A1 => REGISTERS_24_62_port, A2 => n369, B1 => 
                           REGISTERS_26_62_port, B2 => n332, ZN => n2233);
   U2317 : AND4_X1 port map( A1 => n2236, A2 => n2235, A3 => n2234, A4 => n2233
                           , ZN => n2248);
   U2318 : AOI22_X1 port map( A1 => REGISTERS_5_62_port, A2 => n147_port, B1 =>
                           REGISTERS_7_62_port, B2 => n110_port, ZN => n2240);
   U2319 : AOI22_X1 port map( A1 => REGISTERS_1_62_port, A2 => n221, B1 => 
                           REGISTERS_3_62_port, B2 => n184, ZN => n2239);
   U2320 : AOI22_X1 port map( A1 => REGISTERS_4_62_port, A2 => n295, B1 => 
                           REGISTERS_6_62_port, B2 => n258_port, ZN => n2238);
   U2321 : AOI22_X1 port map( A1 => REGISTERS_0_62_port, A2 => n369, B1 => 
                           REGISTERS_2_62_port, B2 => n332, ZN => n2237);
   U2322 : NAND4_X1 port map( A1 => n2240, A2 => n2239, A3 => n2238, A4 => 
                           n2237, ZN => n2246);
   U2323 : AOI22_X1 port map( A1 => REGISTERS_13_62_port, A2 => n147_port, B1 
                           => REGISTERS_15_62_port, B2 => n110_port, ZN => 
                           n2244);
   U2324 : AOI22_X1 port map( A1 => REGISTERS_9_62_port, A2 => n221, B1 => 
                           REGISTERS_11_62_port, B2 => n184, ZN => n2243);
   U2325 : AOI22_X1 port map( A1 => REGISTERS_12_62_port, A2 => n295, B1 => 
                           REGISTERS_14_62_port, B2 => n258_port, ZN => n2242);
   U2326 : AOI22_X1 port map( A1 => REGISTERS_8_62_port, A2 => n369, B1 => 
                           REGISTERS_10_62_port, B2 => n332, ZN => n2241);
   U2327 : NAND4_X1 port map( A1 => n2244, A2 => n2243, A3 => n2242, A4 => 
                           n2241, ZN => n2245);
   U2328 : AOI22_X1 port map( A1 => n2246, A2 => n27, B1 => n2245, B2 => n24, 
                           ZN => n2247);
   U2329 : OAI221_X1 port map( B1 => n2271, B2 => n2249, C1 => n2269, C2 => 
                           n2248, A => n2247, ZN => N97);
   U2330 : AOI22_X1 port map( A1 => REGISTERS_21_63_port, A2 => n148_port, B1 
                           => REGISTERS_23_63_port, B2 => n111_port, ZN => 
                           n2253);
   U2331 : AOI22_X1 port map( A1 => REGISTERS_17_63_port, A2 => n222, B1 => 
                           REGISTERS_19_63_port, B2 => n185, ZN => n2252);
   U2332 : AOI22_X1 port map( A1 => REGISTERS_20_63_port, A2 => n296, B1 => 
                           REGISTERS_22_63_port, B2 => n259_port, ZN => n2251);
   U2333 : AOI22_X1 port map( A1 => REGISTERS_16_63_port, A2 => n370, B1 => 
                           REGISTERS_18_63_port, B2 => n333, ZN => n2250);
   U2334 : AND4_X1 port map( A1 => n2253, A2 => n2252, A3 => n2251, A4 => n2250
                           , ZN => n2272);
   U2335 : AOI22_X1 port map( A1 => REGISTERS_29_63_port, A2 => n148_port, B1 
                           => REGISTERS_31_63_port, B2 => n111_port, ZN => 
                           n2257);
   U2336 : AOI22_X1 port map( A1 => REGISTERS_25_63_port, A2 => n222, B1 => 
                           REGISTERS_27_63_port, B2 => n185, ZN => n2256);
   U2337 : AOI22_X1 port map( A1 => REGISTERS_28_63_port, A2 => n296, B1 => 
                           REGISTERS_30_63_port, B2 => n259_port, ZN => n2255);
   U2338 : AOI22_X1 port map( A1 => REGISTERS_24_63_port, A2 => n370, B1 => 
                           REGISTERS_26_63_port, B2 => n333, ZN => n2254);
   U2339 : AND4_X1 port map( A1 => n2257, A2 => n2256, A3 => n2255, A4 => n2254
                           , ZN => n2270);
   U2340 : AOI22_X1 port map( A1 => REGISTERS_5_63_port, A2 => n148_port, B1 =>
                           REGISTERS_7_63_port, B2 => n111_port, ZN => n2261);
   U2341 : AOI22_X1 port map( A1 => REGISTERS_1_63_port, A2 => n222, B1 => 
                           REGISTERS_3_63_port, B2 => n185, ZN => n2260);
   U2342 : AOI22_X1 port map( A1 => REGISTERS_4_63_port, A2 => n296, B1 => 
                           REGISTERS_6_63_port, B2 => n259_port, ZN => n2259);
   U2343 : AOI22_X1 port map( A1 => REGISTERS_0_63_port, A2 => n370, B1 => 
                           REGISTERS_2_63_port, B2 => n333, ZN => n2258);
   U2344 : NAND4_X1 port map( A1 => n2261, A2 => n2260, A3 => n2259, A4 => 
                           n2258, ZN => n2267);
   U2345 : AOI22_X1 port map( A1 => REGISTERS_13_63_port, A2 => n148_port, B1 
                           => REGISTERS_15_63_port, B2 => n111_port, ZN => 
                           n2265);
   U2346 : AOI22_X1 port map( A1 => REGISTERS_9_63_port, A2 => n222, B1 => 
                           REGISTERS_11_63_port, B2 => n185, ZN => n2264);
   U2347 : AOI22_X1 port map( A1 => REGISTERS_12_63_port, A2 => n296, B1 => 
                           REGISTERS_14_63_port, B2 => n259_port, ZN => n2263);
   U2348 : AOI22_X1 port map( A1 => REGISTERS_8_63_port, A2 => n370, B1 => 
                           REGISTERS_10_63_port, B2 => n333, ZN => n2262);
   U2349 : NAND4_X1 port map( A1 => n2265, A2 => n2264, A3 => n2263, A4 => 
                           n2262, ZN => n2266);
   U2350 : AOI22_X1 port map( A1 => n27, A2 => n2267, B1 => n24, B2 => n2266, 
                           ZN => n2268);
   U2351 : OAI221_X1 port map( B1 => n2272, B2 => n2271, C1 => n2270, C2 => 
                           n2269, A => n2268, ZN => N96);
   U2352 : NOR2_X1 port map( A1 => n5677, A2 => ADD_RD2(1), ZN => n2277);
   U2353 : NOR2_X1 port map( A1 => n5677, A2 => n5676, ZN => n2278);
   U2354 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n423, B1 => 
                           REGISTERS_23_0_port, B2 => n386, ZN => n2284);
   U2355 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n2279);
   U2356 : NOR2_X1 port map( A1 => n5676, A2 => ADD_RD2(2), ZN => n2280);
   U2357 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n497, B1 => 
                           REGISTERS_19_0_port, B2 => n460, ZN => n2283);
   U2358 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n571, B1 => 
                           REGISTERS_22_0_port, B2 => n534, ZN => n2282);
   U2359 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n645, B1 => 
                           REGISTERS_18_0_port, B2 => n608, ZN => n2281);
   U2360 : AND4_X1 port map( A1 => n2284, A2 => n2283, A3 => n2282, A4 => n2281
                           , ZN => n2301);
   U2361 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n423, B1 => 
                           REGISTERS_31_0_port, B2 => n386, ZN => n2288);
   U2362 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n497, B1 => 
                           REGISTERS_27_0_port, B2 => n460, ZN => n2287);
   U2363 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n571, B1 => 
                           REGISTERS_30_0_port, B2 => n534, ZN => n2286);
   U2364 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n645, B1 => 
                           REGISTERS_26_0_port, B2 => n608, ZN => n2285);
   U2365 : AND4_X1 port map( A1 => n2288, A2 => n2287, A3 => n2286, A4 => n2285
                           , ZN => n2300);
   U2366 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n423, B1 => 
                           REGISTERS_7_0_port, B2 => n386, ZN => n2292);
   U2367 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n497, B1 => 
                           REGISTERS_3_0_port, B2 => n460, ZN => n2291);
   U2368 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n571, B1 => 
                           REGISTERS_6_0_port, B2 => n534, ZN => n2290);
   U2369 : AOI22_X1 port map( A1 => REGISTERS_0_0_port, A2 => n645, B1 => 
                           REGISTERS_2_0_port, B2 => n608, ZN => n2289);
   U2370 : NAND4_X1 port map( A1 => n2292, A2 => n2291, A3 => n2290, A4 => 
                           n2289, ZN => n2298);
   U2371 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n423, B1 => 
                           REGISTERS_15_0_port, B2 => n386, ZN => n2296);
   U2372 : AOI22_X1 port map( A1 => REGISTERS_9_0_port, A2 => n497, B1 => 
                           REGISTERS_11_0_port, B2 => n460, ZN => n2295);
   U2373 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n571, B1 => 
                           REGISTERS_14_0_port, B2 => n534, ZN => n2294);
   U2374 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n645, B1 => 
                           REGISTERS_10_0_port, B2 => n608, ZN => n2293);
   U2375 : NAND4_X1 port map( A1 => n2296, A2 => n2295, A3 => n2294, A4 => 
                           n2293, ZN => n2297);
   U2376 : AOI22_X1 port map( A1 => n2298, A2 => n23, B1 => n2297, B2 => n22, 
                           ZN => n2299);
   U2377 : OAI221_X1 port map( B1 => n5673, B2 => n2301, C1 => n5671, C2 => 
                           n2300, A => n2299, ZN => N288);
   U2378 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n423, B1 => 
                           REGISTERS_23_1_port, B2 => n386, ZN => n2305);
   U2379 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n497, B1 => 
                           REGISTERS_19_1_port, B2 => n460, ZN => n2304);
   U2380 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n571, B1 => 
                           REGISTERS_22_1_port, B2 => n534, ZN => n2303);
   U2381 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n645, B1 => 
                           REGISTERS_18_1_port, B2 => n608, ZN => n2302);
   U2382 : AND4_X1 port map( A1 => n2305, A2 => n2304, A3 => n2303, A4 => n2302
                           , ZN => n2322);
   U2383 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n423, B1 => 
                           REGISTERS_31_1_port, B2 => n386, ZN => n2309);
   U2384 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n497, B1 => 
                           REGISTERS_27_1_port, B2 => n460, ZN => n2308);
   U2385 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n571, B1 => 
                           REGISTERS_30_1_port, B2 => n534, ZN => n2307);
   U2386 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n645, B1 => 
                           REGISTERS_26_1_port, B2 => n608, ZN => n2306);
   U2387 : AND4_X1 port map( A1 => n2309, A2 => n2308, A3 => n2307, A4 => n2306
                           , ZN => n2321);
   U2388 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n423, B1 => 
                           REGISTERS_7_1_port, B2 => n386, ZN => n2313);
   U2389 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n497, B1 => 
                           REGISTERS_3_1_port, B2 => n460, ZN => n2312);
   U2390 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n571, B1 => 
                           REGISTERS_6_1_port, B2 => n534, ZN => n2311);
   U2391 : AOI22_X1 port map( A1 => REGISTERS_0_1_port, A2 => n645, B1 => 
                           REGISTERS_2_1_port, B2 => n608, ZN => n2310);
   U2392 : NAND4_X1 port map( A1 => n2313, A2 => n2312, A3 => n2311, A4 => 
                           n2310, ZN => n2319);
   U2393 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n423, B1 => 
                           REGISTERS_15_1_port, B2 => n386, ZN => n2317);
   U2394 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n497, B1 => 
                           REGISTERS_11_1_port, B2 => n460, ZN => n2316);
   U2395 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n571, B1 => 
                           REGISTERS_14_1_port, B2 => n534, ZN => n2315);
   U2396 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n645, B1 => 
                           REGISTERS_10_1_port, B2 => n608, ZN => n2314);
   U2397 : NAND4_X1 port map( A1 => n2317, A2 => n2316, A3 => n2315, A4 => 
                           n2314, ZN => n2318);
   U2398 : AOI22_X1 port map( A1 => n2319, A2 => n23, B1 => n2318, B2 => n22, 
                           ZN => n2320);
   U2399 : OAI221_X1 port map( B1 => n5673, B2 => n2322, C1 => n5671, C2 => 
                           n2321, A => n2320, ZN => N287);
   U2400 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n423, B1 => 
                           REGISTERS_23_2_port, B2 => n386, ZN => n2326);
   U2401 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n497, B1 => 
                           REGISTERS_19_2_port, B2 => n460, ZN => n2325);
   U2402 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n571, B1 => 
                           REGISTERS_22_2_port, B2 => n534, ZN => n2324);
   U2403 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n645, B1 => 
                           REGISTERS_18_2_port, B2 => n608, ZN => n2323);
   U2404 : AND4_X1 port map( A1 => n2326, A2 => n2325, A3 => n2324, A4 => n2323
                           , ZN => n2343);
   U2405 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n423, B1 => 
                           REGISTERS_31_2_port, B2 => n386, ZN => n2330);
   U2406 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n497, B1 => 
                           REGISTERS_27_2_port, B2 => n460, ZN => n2329);
   U2407 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n571, B1 => 
                           REGISTERS_30_2_port, B2 => n534, ZN => n2328);
   U2408 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n645, B1 => 
                           REGISTERS_26_2_port, B2 => n608, ZN => n2327);
   U2409 : AND4_X1 port map( A1 => n2330, A2 => n2329, A3 => n2328, A4 => n2327
                           , ZN => n2342);
   U2410 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n423, B1 => 
                           REGISTERS_7_2_port, B2 => n386, ZN => n2334);
   U2411 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n497, B1 => 
                           REGISTERS_3_2_port, B2 => n460, ZN => n2333);
   U2412 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n571, B1 => 
                           REGISTERS_6_2_port, B2 => n534, ZN => n2332);
   U2413 : AOI22_X1 port map( A1 => REGISTERS_0_2_port, A2 => n645, B1 => 
                           REGISTERS_2_2_port, B2 => n608, ZN => n2331);
   U2414 : NAND4_X1 port map( A1 => n2334, A2 => n2333, A3 => n2332, A4 => 
                           n2331, ZN => n2340);
   U2415 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n423, B1 => 
                           REGISTERS_15_2_port, B2 => n386, ZN => n2338);
   U2416 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n497, B1 => 
                           REGISTERS_11_2_port, B2 => n460, ZN => n2337);
   U2417 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n571, B1 => 
                           REGISTERS_14_2_port, B2 => n534, ZN => n2336);
   U2418 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n645, B1 => 
                           REGISTERS_10_2_port, B2 => n608, ZN => n2335);
   U2419 : NAND4_X1 port map( A1 => n2338, A2 => n2337, A3 => n2336, A4 => 
                           n2335, ZN => n2339);
   U2420 : AOI22_X1 port map( A1 => n2340, A2 => n23, B1 => n2339, B2 => n22, 
                           ZN => n2341);
   U2421 : OAI221_X1 port map( B1 => n5673, B2 => n2343, C1 => n5671, C2 => 
                           n2342, A => n2341, ZN => N286);
   U2422 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n424, B1 => 
                           REGISTERS_23_3_port, B2 => n387, ZN => n2347);
   U2423 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n498, B1 => 
                           REGISTERS_19_3_port, B2 => n461, ZN => n2346);
   U2424 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n572, B1 => 
                           REGISTERS_22_3_port, B2 => n535, ZN => n2345);
   U2425 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n646, B1 => 
                           REGISTERS_18_3_port, B2 => n609, ZN => n2344);
   U2426 : AND4_X1 port map( A1 => n2347, A2 => n2346, A3 => n2345, A4 => n2344
                           , ZN => n2364);
   U2427 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n424, B1 => 
                           REGISTERS_31_3_port, B2 => n387, ZN => n2351);
   U2428 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n498, B1 => 
                           REGISTERS_27_3_port, B2 => n461, ZN => n2350);
   U2429 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n572, B1 => 
                           REGISTERS_30_3_port, B2 => n535, ZN => n2349);
   U2430 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n646, B1 => 
                           REGISTERS_26_3_port, B2 => n609, ZN => n2348);
   U2431 : AND4_X1 port map( A1 => n2351, A2 => n2350, A3 => n2349, A4 => n2348
                           , ZN => n2363);
   U2432 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n424, B1 => 
                           REGISTERS_7_3_port, B2 => n387, ZN => n2355);
   U2433 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n498, B1 => 
                           REGISTERS_3_3_port, B2 => n461, ZN => n2354);
   U2434 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n572, B1 => 
                           REGISTERS_6_3_port, B2 => n535, ZN => n2353);
   U2435 : AOI22_X1 port map( A1 => REGISTERS_0_3_port, A2 => n646, B1 => 
                           REGISTERS_2_3_port, B2 => n609, ZN => n2352);
   U2436 : NAND4_X1 port map( A1 => n2355, A2 => n2354, A3 => n2353, A4 => 
                           n2352, ZN => n2361);
   U2437 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n424, B1 => 
                           REGISTERS_15_3_port, B2 => n387, ZN => n2359);
   U2438 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n498, B1 => 
                           REGISTERS_11_3_port, B2 => n461, ZN => n2358);
   U2439 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n572, B1 => 
                           REGISTERS_14_3_port, B2 => n535, ZN => n2357);
   U2440 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n646, B1 => 
                           REGISTERS_10_3_port, B2 => n609, ZN => n2356);
   U2441 : NAND4_X1 port map( A1 => n2359, A2 => n2358, A3 => n2357, A4 => 
                           n2356, ZN => n2360);
   U2442 : AOI22_X1 port map( A1 => n2361, A2 => n23, B1 => n2360, B2 => n22, 
                           ZN => n2362);
   U2443 : OAI221_X1 port map( B1 => n5673, B2 => n2364, C1 => n5671, C2 => 
                           n2363, A => n2362, ZN => N285);
   U2444 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n424, B1 => 
                           REGISTERS_23_4_port, B2 => n387, ZN => n2368);
   U2445 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n498, B1 => 
                           REGISTERS_19_4_port, B2 => n461, ZN => n2367);
   U2446 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n572, B1 => 
                           REGISTERS_22_4_port, B2 => n535, ZN => n2366);
   U2447 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n646, B1 => 
                           REGISTERS_18_4_port, B2 => n609, ZN => n2365);
   U2448 : AND4_X1 port map( A1 => n2368, A2 => n2367, A3 => n2366, A4 => n2365
                           , ZN => n2385);
   U2449 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n424, B1 => 
                           REGISTERS_31_4_port, B2 => n387, ZN => n2372);
   U2450 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n498, B1 => 
                           REGISTERS_27_4_port, B2 => n461, ZN => n2371);
   U2451 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n572, B1 => 
                           REGISTERS_30_4_port, B2 => n535, ZN => n2370);
   U2452 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n646, B1 => 
                           REGISTERS_26_4_port, B2 => n609, ZN => n2369);
   U2453 : AND4_X1 port map( A1 => n2372, A2 => n2371, A3 => n2370, A4 => n2369
                           , ZN => n2384);
   U2454 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n424, B1 => 
                           REGISTERS_7_4_port, B2 => n387, ZN => n2376);
   U2455 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n498, B1 => 
                           REGISTERS_3_4_port, B2 => n461, ZN => n2375);
   U2456 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n572, B1 => 
                           REGISTERS_6_4_port, B2 => n535, ZN => n2374);
   U2457 : AOI22_X1 port map( A1 => REGISTERS_0_4_port, A2 => n646, B1 => 
                           REGISTERS_2_4_port, B2 => n609, ZN => n2373);
   U2458 : NAND4_X1 port map( A1 => n2376, A2 => n2375, A3 => n2374, A4 => 
                           n2373, ZN => n2382);
   U2459 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n424, B1 => 
                           REGISTERS_15_4_port, B2 => n387, ZN => n2380);
   U2460 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n498, B1 => 
                           REGISTERS_11_4_port, B2 => n461, ZN => n2379);
   U2461 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n572, B1 => 
                           REGISTERS_14_4_port, B2 => n535, ZN => n2378);
   U2462 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n646, B1 => 
                           REGISTERS_10_4_port, B2 => n609, ZN => n2377);
   U2463 : NAND4_X1 port map( A1 => n2380, A2 => n2379, A3 => n2378, A4 => 
                           n2377, ZN => n2381);
   U2464 : AOI22_X1 port map( A1 => n2382, A2 => n23, B1 => n2381, B2 => n22, 
                           ZN => n2383);
   U2465 : OAI221_X1 port map( B1 => n5673, B2 => n2385, C1 => n5671, C2 => 
                           n2384, A => n2383, ZN => N284);
   U2466 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n424, B1 => 
                           REGISTERS_23_5_port, B2 => n387, ZN => n2389);
   U2467 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n498, B1 => 
                           REGISTERS_19_5_port, B2 => n461, ZN => n2388);
   U2468 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n572, B1 => 
                           REGISTERS_22_5_port, B2 => n535, ZN => n2387);
   U2469 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n646, B1 => 
                           REGISTERS_18_5_port, B2 => n609, ZN => n2386);
   U2470 : AND4_X1 port map( A1 => n2389, A2 => n2388, A3 => n2387, A4 => n2386
                           , ZN => n2406);
   U2471 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n424, B1 => 
                           REGISTERS_31_5_port, B2 => n387, ZN => n2393);
   U2472 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n498, B1 => 
                           REGISTERS_27_5_port, B2 => n461, ZN => n2392);
   U2473 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n572, B1 => 
                           REGISTERS_30_5_port, B2 => n535, ZN => n2391);
   U2474 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n646, B1 => 
                           REGISTERS_26_5_port, B2 => n609, ZN => n2390);
   U2475 : AND4_X1 port map( A1 => n2393, A2 => n2392, A3 => n2391, A4 => n2390
                           , ZN => n2405);
   U2476 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n424, B1 => 
                           REGISTERS_7_5_port, B2 => n387, ZN => n2397);
   U2477 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n498, B1 => 
                           REGISTERS_3_5_port, B2 => n461, ZN => n2396);
   U2478 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n572, B1 => 
                           REGISTERS_6_5_port, B2 => n535, ZN => n2395);
   U2479 : AOI22_X1 port map( A1 => REGISTERS_0_5_port, A2 => n646, B1 => 
                           REGISTERS_2_5_port, B2 => n609, ZN => n2394);
   U2480 : NAND4_X1 port map( A1 => n2397, A2 => n2396, A3 => n2395, A4 => 
                           n2394, ZN => n2403);
   U2481 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n424, B1 => 
                           REGISTERS_15_5_port, B2 => n387, ZN => n2401);
   U2482 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n498, B1 => 
                           REGISTERS_11_5_port, B2 => n461, ZN => n2400);
   U2483 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n572, B1 => 
                           REGISTERS_14_5_port, B2 => n535, ZN => n2399);
   U2484 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n646, B1 => 
                           REGISTERS_10_5_port, B2 => n609, ZN => n2398);
   U2485 : NAND4_X1 port map( A1 => n2401, A2 => n2400, A3 => n2399, A4 => 
                           n2398, ZN => n2402);
   U2486 : AOI22_X1 port map( A1 => n2403, A2 => n23, B1 => n2402, B2 => n22, 
                           ZN => n2404);
   U2487 : OAI221_X1 port map( B1 => n5673, B2 => n2406, C1 => n5671, C2 => 
                           n2405, A => n2404, ZN => N283);
   U2488 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n425, B1 => 
                           REGISTERS_23_6_port, B2 => n388, ZN => n2410);
   U2489 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n499, B1 => 
                           REGISTERS_19_6_port, B2 => n462, ZN => n2409);
   U2490 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n573, B1 => 
                           REGISTERS_22_6_port, B2 => n536, ZN => n2408);
   U2491 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n647, B1 => 
                           REGISTERS_18_6_port, B2 => n610, ZN => n2407);
   U2492 : AND4_X1 port map( A1 => n2410, A2 => n2409, A3 => n2408, A4 => n2407
                           , ZN => n2427);
   U2493 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n425, B1 => 
                           REGISTERS_31_6_port, B2 => n388, ZN => n2414);
   U2494 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n499, B1 => 
                           REGISTERS_27_6_port, B2 => n462, ZN => n2413);
   U2495 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n573, B1 => 
                           REGISTERS_30_6_port, B2 => n536, ZN => n2412);
   U2496 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n647, B1 => 
                           REGISTERS_26_6_port, B2 => n610, ZN => n2411);
   U2497 : AND4_X1 port map( A1 => n2414, A2 => n2413, A3 => n2412, A4 => n2411
                           , ZN => n2426);
   U2498 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n425, B1 => 
                           REGISTERS_7_6_port, B2 => n388, ZN => n2418);
   U2499 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n499, B1 => 
                           REGISTERS_3_6_port, B2 => n462, ZN => n2417);
   U2500 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n573, B1 => 
                           REGISTERS_6_6_port, B2 => n536, ZN => n2416);
   U2501 : AOI22_X1 port map( A1 => REGISTERS_0_6_port, A2 => n647, B1 => 
                           REGISTERS_2_6_port, B2 => n610, ZN => n2415);
   U2502 : NAND4_X1 port map( A1 => n2418, A2 => n2417, A3 => n2416, A4 => 
                           n2415, ZN => n2424);
   U2503 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n425, B1 => 
                           REGISTERS_15_6_port, B2 => n388, ZN => n2422);
   U2504 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n499, B1 => 
                           REGISTERS_11_6_port, B2 => n462, ZN => n2421);
   U2505 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n573, B1 => 
                           REGISTERS_14_6_port, B2 => n536, ZN => n2420);
   U2506 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n647, B1 => 
                           REGISTERS_10_6_port, B2 => n610, ZN => n2419);
   U2507 : NAND4_X1 port map( A1 => n2422, A2 => n2421, A3 => n2420, A4 => 
                           n2419, ZN => n2423);
   U2508 : AOI22_X1 port map( A1 => n2424, A2 => n23, B1 => n2423, B2 => n22, 
                           ZN => n2425);
   U2509 : OAI221_X1 port map( B1 => n5673, B2 => n2427, C1 => n5671, C2 => 
                           n2426, A => n2425, ZN => N282);
   U2510 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n425, B1 => 
                           REGISTERS_23_7_port, B2 => n388, ZN => n2431);
   U2511 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n499, B1 => 
                           REGISTERS_19_7_port, B2 => n462, ZN => n2430);
   U2512 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n573, B1 => 
                           REGISTERS_22_7_port, B2 => n536, ZN => n2429);
   U2513 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n647, B1 => 
                           REGISTERS_18_7_port, B2 => n610, ZN => n2428);
   U2514 : AND4_X1 port map( A1 => n2431, A2 => n2430, A3 => n2429, A4 => n2428
                           , ZN => n2448);
   U2515 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n425, B1 => 
                           REGISTERS_31_7_port, B2 => n388, ZN => n2435);
   U2516 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n499, B1 => 
                           REGISTERS_27_7_port, B2 => n462, ZN => n2434);
   U2517 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n573, B1 => 
                           REGISTERS_30_7_port, B2 => n536, ZN => n2433);
   U2518 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n647, B1 => 
                           REGISTERS_26_7_port, B2 => n610, ZN => n2432);
   U2519 : AND4_X1 port map( A1 => n2435, A2 => n2434, A3 => n2433, A4 => n2432
                           , ZN => n2447);
   U2520 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n425, B1 => 
                           REGISTERS_7_7_port, B2 => n388, ZN => n2439);
   U2521 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n499, B1 => 
                           REGISTERS_3_7_port, B2 => n462, ZN => n2438);
   U2522 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n573, B1 => 
                           REGISTERS_6_7_port, B2 => n536, ZN => n2437);
   U2523 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n647, B1 => 
                           REGISTERS_2_7_port, B2 => n610, ZN => n2436);
   U2524 : NAND4_X1 port map( A1 => n2439, A2 => n2438, A3 => n2437, A4 => 
                           n2436, ZN => n2445);
   U2525 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n425, B1 => 
                           REGISTERS_15_7_port, B2 => n388, ZN => n2443);
   U2526 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n499, B1 => 
                           REGISTERS_11_7_port, B2 => n462, ZN => n2442);
   U2527 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n573, B1 => 
                           REGISTERS_14_7_port, B2 => n536, ZN => n2441);
   U2528 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n647, B1 => 
                           REGISTERS_10_7_port, B2 => n610, ZN => n2440);
   U2529 : NAND4_X1 port map( A1 => n2443, A2 => n2442, A3 => n2441, A4 => 
                           n2440, ZN => n2444);
   U2530 : AOI22_X1 port map( A1 => n2445, A2 => n23, B1 => n2444, B2 => n22, 
                           ZN => n2446);
   U2531 : OAI221_X1 port map( B1 => n5673, B2 => n2448, C1 => n5671, C2 => 
                           n2447, A => n2446, ZN => N281);
   U2532 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n425, B1 => 
                           REGISTERS_23_8_port, B2 => n388, ZN => n2452);
   U2533 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n499, B1 => 
                           REGISTERS_19_8_port, B2 => n462, ZN => n2451);
   U2534 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n573, B1 => 
                           REGISTERS_22_8_port, B2 => n536, ZN => n2450);
   U2535 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n647, B1 => 
                           REGISTERS_18_8_port, B2 => n610, ZN => n2449);
   U2536 : AND4_X1 port map( A1 => n2452, A2 => n2451, A3 => n2450, A4 => n2449
                           , ZN => n4517);
   U2537 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n425, B1 => 
                           REGISTERS_31_8_port, B2 => n388, ZN => n4504);
   U2538 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n499, B1 => 
                           REGISTERS_27_8_port, B2 => n462, ZN => n2455);
   U2539 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n573, B1 => 
                           REGISTERS_30_8_port, B2 => n536, ZN => n2454);
   U2540 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n647, B1 => 
                           REGISTERS_26_8_port, B2 => n610, ZN => n2453);
   U2541 : AND4_X1 port map( A1 => n4504, A2 => n2455, A3 => n2454, A4 => n2453
                           , ZN => n4516);
   U2542 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n425, B1 => 
                           REGISTERS_7_8_port, B2 => n388, ZN => n4508);
   U2543 : AOI22_X1 port map( A1 => REGISTERS_1_8_port, A2 => n499, B1 => 
                           REGISTERS_3_8_port, B2 => n462, ZN => n4507);
   U2544 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n573, B1 => 
                           REGISTERS_6_8_port, B2 => n536, ZN => n4506);
   U2545 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n647, B1 => 
                           REGISTERS_2_8_port, B2 => n610, ZN => n4505);
   U2546 : NAND4_X1 port map( A1 => n4508, A2 => n4507, A3 => n4506, A4 => 
                           n4505, ZN => n4514);
   U2547 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n425, B1 => 
                           REGISTERS_15_8_port, B2 => n388, ZN => n4512);
   U2548 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n499, B1 => 
                           REGISTERS_11_8_port, B2 => n462, ZN => n4511);
   U2549 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n573, B1 => 
                           REGISTERS_14_8_port, B2 => n536, ZN => n4510);
   U2550 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n647, B1 => 
                           REGISTERS_10_8_port, B2 => n610, ZN => n4509);
   U2551 : NAND4_X1 port map( A1 => n4512, A2 => n4511, A3 => n4510, A4 => 
                           n4509, ZN => n4513);
   U2552 : AOI22_X1 port map( A1 => n4514, A2 => n23, B1 => n4513, B2 => n22, 
                           ZN => n4515);
   U2553 : OAI221_X1 port map( B1 => n5673, B2 => n4517, C1 => n5671, C2 => 
                           n4516, A => n4515, ZN => N280);
   U2554 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n426, B1 => 
                           REGISTERS_23_9_port, B2 => n389, ZN => n4521);
   U2555 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n500, B1 => 
                           REGISTERS_19_9_port, B2 => n463, ZN => n4520);
   U2556 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n574, B1 => 
                           REGISTERS_22_9_port, B2 => n537, ZN => n4519);
   U2557 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n648, B1 => 
                           REGISTERS_18_9_port, B2 => n611, ZN => n4518);
   U2558 : AND4_X1 port map( A1 => n4521, A2 => n4520, A3 => n4519, A4 => n4518
                           , ZN => n4538);
   U2559 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n426, B1 => 
                           REGISTERS_31_9_port, B2 => n389, ZN => n4525);
   U2560 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n500, B1 => 
                           REGISTERS_27_9_port, B2 => n463, ZN => n4524);
   U2561 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n574, B1 => 
                           REGISTERS_30_9_port, B2 => n537, ZN => n4523);
   U2562 : AOI22_X1 port map( A1 => REGISTERS_24_9_port, A2 => n648, B1 => 
                           REGISTERS_26_9_port, B2 => n611, ZN => n4522);
   U2563 : AND4_X1 port map( A1 => n4525, A2 => n4524, A3 => n4523, A4 => n4522
                           , ZN => n4537);
   U2564 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n426, B1 => 
                           REGISTERS_7_9_port, B2 => n389, ZN => n4529);
   U2565 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n500, B1 => 
                           REGISTERS_3_9_port, B2 => n463, ZN => n4528);
   U2566 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n574, B1 => 
                           REGISTERS_6_9_port, B2 => n537, ZN => n4527);
   U2567 : AOI22_X1 port map( A1 => REGISTERS_0_9_port, A2 => n648, B1 => 
                           REGISTERS_2_9_port, B2 => n611, ZN => n4526);
   U2568 : NAND4_X1 port map( A1 => n4529, A2 => n4528, A3 => n4527, A4 => 
                           n4526, ZN => n4535);
   U2569 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n426, B1 => 
                           REGISTERS_15_9_port, B2 => n389, ZN => n4533);
   U2570 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n500, B1 => 
                           REGISTERS_11_9_port, B2 => n463, ZN => n4532);
   U2571 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n574, B1 => 
                           REGISTERS_14_9_port, B2 => n537, ZN => n4531);
   U2572 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n648, B1 => 
                           REGISTERS_10_9_port, B2 => n611, ZN => n4530);
   U2573 : NAND4_X1 port map( A1 => n4533, A2 => n4532, A3 => n4531, A4 => 
                           n4530, ZN => n4534);
   U2574 : AOI22_X1 port map( A1 => n4535, A2 => n23, B1 => n4534, B2 => n22, 
                           ZN => n4536);
   U2575 : OAI221_X1 port map( B1 => n5673, B2 => n4538, C1 => n5671, C2 => 
                           n4537, A => n4536, ZN => N279);
   U2576 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n426, B1 => 
                           REGISTERS_23_10_port, B2 => n389, ZN => n4542);
   U2577 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n500, B1 => 
                           REGISTERS_19_10_port, B2 => n463, ZN => n4541);
   U2578 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n574, B1 => 
                           REGISTERS_22_10_port, B2 => n537, ZN => n4540);
   U2579 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n648, B1 => 
                           REGISTERS_18_10_port, B2 => n611, ZN => n4539);
   U2580 : AND4_X1 port map( A1 => n4542, A2 => n4541, A3 => n4540, A4 => n4539
                           , ZN => n4559);
   U2581 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n426, B1 => 
                           REGISTERS_31_10_port, B2 => n389, ZN => n4546);
   U2582 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n500, B1 => 
                           REGISTERS_27_10_port, B2 => n463, ZN => n4545);
   U2583 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n574, B1 => 
                           REGISTERS_30_10_port, B2 => n537, ZN => n4544);
   U2584 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n648, B1 => 
                           REGISTERS_26_10_port, B2 => n611, ZN => n4543);
   U2585 : AND4_X1 port map( A1 => n4546, A2 => n4545, A3 => n4544, A4 => n4543
                           , ZN => n4558);
   U2586 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n426, B1 => 
                           REGISTERS_7_10_port, B2 => n389, ZN => n4550);
   U2587 : AOI22_X1 port map( A1 => REGISTERS_1_10_port, A2 => n500, B1 => 
                           REGISTERS_3_10_port, B2 => n463, ZN => n4549);
   U2588 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n574, B1 => 
                           REGISTERS_6_10_port, B2 => n537, ZN => n4548);
   U2589 : AOI22_X1 port map( A1 => REGISTERS_0_10_port, A2 => n648, B1 => 
                           REGISTERS_2_10_port, B2 => n611, ZN => n4547);
   U2590 : NAND4_X1 port map( A1 => n4550, A2 => n4549, A3 => n4548, A4 => 
                           n4547, ZN => n4556);
   U2591 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n426, B1 => 
                           REGISTERS_15_10_port, B2 => n389, ZN => n4554);
   U2592 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n500, B1 => 
                           REGISTERS_11_10_port, B2 => n463, ZN => n4553);
   U2593 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n574, B1 => 
                           REGISTERS_14_10_port, B2 => n537, ZN => n4552);
   U2594 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n648, B1 => 
                           REGISTERS_10_10_port, B2 => n611, ZN => n4551);
   U2595 : NAND4_X1 port map( A1 => n4554, A2 => n4553, A3 => n4552, A4 => 
                           n4551, ZN => n4555);
   U2596 : AOI22_X1 port map( A1 => n4556, A2 => n23, B1 => n4555, B2 => n22, 
                           ZN => n4557);
   U2597 : OAI221_X1 port map( B1 => n5673, B2 => n4559, C1 => n5671, C2 => 
                           n4558, A => n4557, ZN => N278);
   U2598 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n426, B1 => 
                           REGISTERS_23_11_port, B2 => n389, ZN => n4563);
   U2599 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n500, B1 => 
                           REGISTERS_19_11_port, B2 => n463, ZN => n4562);
   U2600 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n574, B1 => 
                           REGISTERS_22_11_port, B2 => n537, ZN => n4561);
   U2601 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n648, B1 => 
                           REGISTERS_18_11_port, B2 => n611, ZN => n4560);
   U2602 : AND4_X1 port map( A1 => n4563, A2 => n4562, A3 => n4561, A4 => n4560
                           , ZN => n4580);
   U2603 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n426, B1 => 
                           REGISTERS_31_11_port, B2 => n389, ZN => n4567);
   U2604 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n500, B1 => 
                           REGISTERS_27_11_port, B2 => n463, ZN => n4566);
   U2605 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n574, B1 => 
                           REGISTERS_30_11_port, B2 => n537, ZN => n4565);
   U2606 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n648, B1 => 
                           REGISTERS_26_11_port, B2 => n611, ZN => n4564);
   U2607 : AND4_X1 port map( A1 => n4567, A2 => n4566, A3 => n4565, A4 => n4564
                           , ZN => n4579);
   U2608 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n426, B1 => 
                           REGISTERS_7_11_port, B2 => n389, ZN => n4571);
   U2609 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n500, B1 => 
                           REGISTERS_3_11_port, B2 => n463, ZN => n4570);
   U2610 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n574, B1 => 
                           REGISTERS_6_11_port, B2 => n537, ZN => n4569);
   U2611 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n648, B1 => 
                           REGISTERS_2_11_port, B2 => n611, ZN => n4568);
   U2612 : NAND4_X1 port map( A1 => n4571, A2 => n4570, A3 => n4569, A4 => 
                           n4568, ZN => n4577);
   U2613 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n426, B1 => 
                           REGISTERS_15_11_port, B2 => n389, ZN => n4575);
   U2614 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n500, B1 => 
                           REGISTERS_11_11_port, B2 => n463, ZN => n4574);
   U2615 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n574, B1 => 
                           REGISTERS_14_11_port, B2 => n537, ZN => n4573);
   U2616 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n648, B1 => 
                           REGISTERS_10_11_port, B2 => n611, ZN => n4572);
   U2617 : NAND4_X1 port map( A1 => n4575, A2 => n4574, A3 => n4573, A4 => 
                           n4572, ZN => n4576);
   U2618 : AOI22_X1 port map( A1 => n4577, A2 => n23, B1 => n4576, B2 => n22, 
                           ZN => n4578);
   U2619 : OAI221_X1 port map( B1 => n5673, B2 => n4580, C1 => n5671, C2 => 
                           n4579, A => n4578, ZN => N277);
   U2620 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n427, B1 => 
                           REGISTERS_23_12_port, B2 => n390, ZN => n4584);
   U2621 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n501, B1 => 
                           REGISTERS_19_12_port, B2 => n464, ZN => n4583);
   U2622 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n575, B1 => 
                           REGISTERS_22_12_port, B2 => n538, ZN => n4582);
   U2623 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n649, B1 => 
                           REGISTERS_18_12_port, B2 => n612, ZN => n4581);
   U2624 : AND4_X1 port map( A1 => n4584, A2 => n4583, A3 => n4582, A4 => n4581
                           , ZN => n4601);
   U2625 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n427, B1 => 
                           REGISTERS_31_12_port, B2 => n390, ZN => n4588);
   U2626 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n501, B1 => 
                           REGISTERS_27_12_port, B2 => n464, ZN => n4587);
   U2627 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n575, B1 => 
                           REGISTERS_30_12_port, B2 => n538, ZN => n4586);
   U2628 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n649, B1 => 
                           REGISTERS_26_12_port, B2 => n612, ZN => n4585);
   U2629 : AND4_X1 port map( A1 => n4588, A2 => n4587, A3 => n4586, A4 => n4585
                           , ZN => n4600);
   U2630 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n427, B1 => 
                           REGISTERS_7_12_port, B2 => n390, ZN => n4592);
   U2631 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n501, B1 => 
                           REGISTERS_3_12_port, B2 => n464, ZN => n4591);
   U2632 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n575, B1 => 
                           REGISTERS_6_12_port, B2 => n538, ZN => n4590);
   U2633 : AOI22_X1 port map( A1 => REGISTERS_0_12_port, A2 => n649, B1 => 
                           REGISTERS_2_12_port, B2 => n612, ZN => n4589);
   U2634 : NAND4_X1 port map( A1 => n4592, A2 => n4591, A3 => n4590, A4 => 
                           n4589, ZN => n4598);
   U2635 : AOI22_X1 port map( A1 => REGISTERS_13_12_port, A2 => n427, B1 => 
                           REGISTERS_15_12_port, B2 => n390, ZN => n4596);
   U2636 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n501, B1 => 
                           REGISTERS_11_12_port, B2 => n464, ZN => n4595);
   U2637 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n575, B1 => 
                           REGISTERS_14_12_port, B2 => n538, ZN => n4594);
   U2638 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n649, B1 => 
                           REGISTERS_10_12_port, B2 => n612, ZN => n4593);
   U2639 : NAND4_X1 port map( A1 => n4596, A2 => n4595, A3 => n4594, A4 => 
                           n4593, ZN => n4597);
   U2640 : AOI22_X1 port map( A1 => n4598, A2 => n23, B1 => n4597, B2 => n22, 
                           ZN => n4599);
   U2641 : OAI221_X1 port map( B1 => n5673, B2 => n4601, C1 => n5671, C2 => 
                           n4600, A => n4599, ZN => N276);
   U2642 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n427, B1 => 
                           REGISTERS_23_13_port, B2 => n390, ZN => n4605);
   U2643 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n501, B1 => 
                           REGISTERS_19_13_port, B2 => n464, ZN => n4604);
   U2644 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n575, B1 => 
                           REGISTERS_22_13_port, B2 => n538, ZN => n4603);
   U2645 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n649, B1 => 
                           REGISTERS_18_13_port, B2 => n612, ZN => n4602);
   U2646 : AND4_X1 port map( A1 => n4605, A2 => n4604, A3 => n4603, A4 => n4602
                           , ZN => n4622);
   U2647 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n427, B1 => 
                           REGISTERS_31_13_port, B2 => n390, ZN => n4609);
   U2648 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n501, B1 => 
                           REGISTERS_27_13_port, B2 => n464, ZN => n4608);
   U2649 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n575, B1 => 
                           REGISTERS_30_13_port, B2 => n538, ZN => n4607);
   U2650 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n649, B1 => 
                           REGISTERS_26_13_port, B2 => n612, ZN => n4606);
   U2651 : AND4_X1 port map( A1 => n4609, A2 => n4608, A3 => n4607, A4 => n4606
                           , ZN => n4621);
   U2652 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n427, B1 => 
                           REGISTERS_7_13_port, B2 => n390, ZN => n4613);
   U2653 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n501, B1 => 
                           REGISTERS_3_13_port, B2 => n464, ZN => n4612);
   U2654 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n575, B1 => 
                           REGISTERS_6_13_port, B2 => n538, ZN => n4611);
   U2655 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n649, B1 => 
                           REGISTERS_2_13_port, B2 => n612, ZN => n4610);
   U2656 : NAND4_X1 port map( A1 => n4613, A2 => n4612, A3 => n4611, A4 => 
                           n4610, ZN => n4619);
   U2657 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n427, B1 => 
                           REGISTERS_15_13_port, B2 => n390, ZN => n4617);
   U2658 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n501, B1 => 
                           REGISTERS_11_13_port, B2 => n464, ZN => n4616);
   U2659 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n575, B1 => 
                           REGISTERS_14_13_port, B2 => n538, ZN => n4615);
   U2660 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n649, B1 => 
                           REGISTERS_10_13_port, B2 => n612, ZN => n4614);
   U2661 : NAND4_X1 port map( A1 => n4617, A2 => n4616, A3 => n4615, A4 => 
                           n4614, ZN => n4618);
   U2662 : AOI22_X1 port map( A1 => n4619, A2 => n23, B1 => n4618, B2 => n22, 
                           ZN => n4620);
   U2663 : OAI221_X1 port map( B1 => n5673, B2 => n4622, C1 => n5671, C2 => 
                           n4621, A => n4620, ZN => N275);
   U2664 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n427, B1 => 
                           REGISTERS_23_14_port, B2 => n390, ZN => n4626);
   U2665 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n501, B1 => 
                           REGISTERS_19_14_port, B2 => n464, ZN => n4625);
   U2666 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n575, B1 => 
                           REGISTERS_22_14_port, B2 => n538, ZN => n4624);
   U2667 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n649, B1 => 
                           REGISTERS_18_14_port, B2 => n612, ZN => n4623);
   U2668 : AND4_X1 port map( A1 => n4626, A2 => n4625, A3 => n4624, A4 => n4623
                           , ZN => n4643);
   U2669 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n427, B1 => 
                           REGISTERS_31_14_port, B2 => n390, ZN => n4630);
   U2670 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n501, B1 => 
                           REGISTERS_27_14_port, B2 => n464, ZN => n4629);
   U2671 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n575, B1 => 
                           REGISTERS_30_14_port, B2 => n538, ZN => n4628);
   U2672 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n649, B1 => 
                           REGISTERS_26_14_port, B2 => n612, ZN => n4627);
   U2673 : AND4_X1 port map( A1 => n4630, A2 => n4629, A3 => n4628, A4 => n4627
                           , ZN => n4642);
   U2674 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n427, B1 => 
                           REGISTERS_7_14_port, B2 => n390, ZN => n4634);
   U2675 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n501, B1 => 
                           REGISTERS_3_14_port, B2 => n464, ZN => n4633);
   U2676 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n575, B1 => 
                           REGISTERS_6_14_port, B2 => n538, ZN => n4632);
   U2677 : AOI22_X1 port map( A1 => REGISTERS_0_14_port, A2 => n649, B1 => 
                           REGISTERS_2_14_port, B2 => n612, ZN => n4631);
   U2678 : NAND4_X1 port map( A1 => n4634, A2 => n4633, A3 => n4632, A4 => 
                           n4631, ZN => n4640);
   U2679 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n427, B1 => 
                           REGISTERS_15_14_port, B2 => n390, ZN => n4638);
   U2680 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n501, B1 => 
                           REGISTERS_11_14_port, B2 => n464, ZN => n4637);
   U2681 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n575, B1 => 
                           REGISTERS_14_14_port, B2 => n538, ZN => n4636);
   U2682 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n649, B1 => 
                           REGISTERS_10_14_port, B2 => n612, ZN => n4635);
   U2683 : NAND4_X1 port map( A1 => n4638, A2 => n4637, A3 => n4636, A4 => 
                           n4635, ZN => n4639);
   U2684 : AOI22_X1 port map( A1 => n4640, A2 => n23, B1 => n4639, B2 => n22, 
                           ZN => n4641);
   U2685 : OAI221_X1 port map( B1 => n5673, B2 => n4643, C1 => n5671, C2 => 
                           n4642, A => n4641, ZN => N274);
   U2686 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n428, B1 => 
                           REGISTERS_23_15_port, B2 => n391, ZN => n4647);
   U2687 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n502, B1 => 
                           REGISTERS_19_15_port, B2 => n465, ZN => n4646);
   U2688 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n576, B1 => 
                           REGISTERS_22_15_port, B2 => n539, ZN => n4645);
   U2689 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n650, B1 => 
                           REGISTERS_18_15_port, B2 => n613, ZN => n4644);
   U2690 : AND4_X1 port map( A1 => n4647, A2 => n4646, A3 => n4645, A4 => n4644
                           , ZN => n4664);
   U2691 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n428, B1 => 
                           REGISTERS_31_15_port, B2 => n391, ZN => n4651);
   U2692 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n502, B1 => 
                           REGISTERS_27_15_port, B2 => n465, ZN => n4650);
   U2693 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n576, B1 => 
                           REGISTERS_30_15_port, B2 => n539, ZN => n4649);
   U2694 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n650, B1 => 
                           REGISTERS_26_15_port, B2 => n613, ZN => n4648);
   U2695 : AND4_X1 port map( A1 => n4651, A2 => n4650, A3 => n4649, A4 => n4648
                           , ZN => n4663);
   U2696 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n428, B1 => 
                           REGISTERS_7_15_port, B2 => n391, ZN => n4655);
   U2697 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n502, B1 => 
                           REGISTERS_3_15_port, B2 => n465, ZN => n4654);
   U2698 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n576, B1 => 
                           REGISTERS_6_15_port, B2 => n539, ZN => n4653);
   U2699 : AOI22_X1 port map( A1 => REGISTERS_0_15_port, A2 => n650, B1 => 
                           REGISTERS_2_15_port, B2 => n613, ZN => n4652);
   U2700 : NAND4_X1 port map( A1 => n4655, A2 => n4654, A3 => n4653, A4 => 
                           n4652, ZN => n4661);
   U2701 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n428, B1 => 
                           REGISTERS_15_15_port, B2 => n391, ZN => n4659);
   U2702 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n502, B1 => 
                           REGISTERS_11_15_port, B2 => n465, ZN => n4658);
   U2703 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n576, B1 => 
                           REGISTERS_14_15_port, B2 => n539, ZN => n4657);
   U2704 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n650, B1 => 
                           REGISTERS_10_15_port, B2 => n613, ZN => n4656);
   U2705 : NAND4_X1 port map( A1 => n4659, A2 => n4658, A3 => n4657, A4 => 
                           n4656, ZN => n4660);
   U2706 : AOI22_X1 port map( A1 => n4661, A2 => n23, B1 => n4660, B2 => n22, 
                           ZN => n4662);
   U2707 : OAI221_X1 port map( B1 => n5673, B2 => n4664, C1 => n5671, C2 => 
                           n4663, A => n4662, ZN => N273);
   U2708 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n428, B1 => 
                           REGISTERS_23_16_port, B2 => n391, ZN => n4668);
   U2709 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n502, B1 => 
                           REGISTERS_19_16_port, B2 => n465, ZN => n4667);
   U2710 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n576, B1 => 
                           REGISTERS_22_16_port, B2 => n539, ZN => n4666);
   U2711 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n650, B1 => 
                           REGISTERS_18_16_port, B2 => n613, ZN => n4665);
   U2712 : AND4_X1 port map( A1 => n4668, A2 => n4667, A3 => n4666, A4 => n4665
                           , ZN => n4685);
   U2713 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n428, B1 => 
                           REGISTERS_31_16_port, B2 => n391, ZN => n4672);
   U2714 : AOI22_X1 port map( A1 => REGISTERS_25_16_port, A2 => n502, B1 => 
                           REGISTERS_27_16_port, B2 => n465, ZN => n4671);
   U2715 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n576, B1 => 
                           REGISTERS_30_16_port, B2 => n539, ZN => n4670);
   U2716 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n650, B1 => 
                           REGISTERS_26_16_port, B2 => n613, ZN => n4669);
   U2717 : AND4_X1 port map( A1 => n4672, A2 => n4671, A3 => n4670, A4 => n4669
                           , ZN => n4684);
   U2718 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n428, B1 => 
                           REGISTERS_7_16_port, B2 => n391, ZN => n4676);
   U2719 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n502, B1 => 
                           REGISTERS_3_16_port, B2 => n465, ZN => n4675);
   U2720 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n576, B1 => 
                           REGISTERS_6_16_port, B2 => n539, ZN => n4674);
   U2721 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n650, B1 => 
                           REGISTERS_2_16_port, B2 => n613, ZN => n4673);
   U2722 : NAND4_X1 port map( A1 => n4676, A2 => n4675, A3 => n4674, A4 => 
                           n4673, ZN => n4682);
   U2723 : AOI22_X1 port map( A1 => REGISTERS_13_16_port, A2 => n428, B1 => 
                           REGISTERS_15_16_port, B2 => n391, ZN => n4680);
   U2724 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n502, B1 => 
                           REGISTERS_11_16_port, B2 => n465, ZN => n4679);
   U2725 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n576, B1 => 
                           REGISTERS_14_16_port, B2 => n539, ZN => n4678);
   U2726 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n650, B1 => 
                           REGISTERS_10_16_port, B2 => n613, ZN => n4677);
   U2727 : NAND4_X1 port map( A1 => n4680, A2 => n4679, A3 => n4678, A4 => 
                           n4677, ZN => n4681);
   U2728 : AOI22_X1 port map( A1 => n4682, A2 => n23, B1 => n4681, B2 => n22, 
                           ZN => n4683);
   U2729 : OAI221_X1 port map( B1 => n5673, B2 => n4685, C1 => n5671, C2 => 
                           n4684, A => n4683, ZN => N272);
   U2730 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n428, B1 => 
                           REGISTERS_23_17_port, B2 => n391, ZN => n4689);
   U2731 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n502, B1 => 
                           REGISTERS_19_17_port, B2 => n465, ZN => n4688);
   U2732 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n576, B1 => 
                           REGISTERS_22_17_port, B2 => n539, ZN => n4687);
   U2733 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n650, B1 => 
                           REGISTERS_18_17_port, B2 => n613, ZN => n4686);
   U2734 : AND4_X1 port map( A1 => n4689, A2 => n4688, A3 => n4687, A4 => n4686
                           , ZN => n4706);
   U2735 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n428, B1 => 
                           REGISTERS_31_17_port, B2 => n391, ZN => n4693);
   U2736 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n502, B1 => 
                           REGISTERS_27_17_port, B2 => n465, ZN => n4692);
   U2737 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n576, B1 => 
                           REGISTERS_30_17_port, B2 => n539, ZN => n4691);
   U2738 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n650, B1 => 
                           REGISTERS_26_17_port, B2 => n613, ZN => n4690);
   U2739 : AND4_X1 port map( A1 => n4693, A2 => n4692, A3 => n4691, A4 => n4690
                           , ZN => n4705);
   U2740 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n428, B1 => 
                           REGISTERS_7_17_port, B2 => n391, ZN => n4697);
   U2741 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n502, B1 => 
                           REGISTERS_3_17_port, B2 => n465, ZN => n4696);
   U2742 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n576, B1 => 
                           REGISTERS_6_17_port, B2 => n539, ZN => n4695);
   U2743 : AOI22_X1 port map( A1 => REGISTERS_0_17_port, A2 => n650, B1 => 
                           REGISTERS_2_17_port, B2 => n613, ZN => n4694);
   U2744 : NAND4_X1 port map( A1 => n4697, A2 => n4696, A3 => n4695, A4 => 
                           n4694, ZN => n4703);
   U2745 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n428, B1 => 
                           REGISTERS_15_17_port, B2 => n391, ZN => n4701);
   U2746 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n502, B1 => 
                           REGISTERS_11_17_port, B2 => n465, ZN => n4700);
   U2747 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n576, B1 => 
                           REGISTERS_14_17_port, B2 => n539, ZN => n4699);
   U2748 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n650, B1 => 
                           REGISTERS_10_17_port, B2 => n613, ZN => n4698);
   U2749 : NAND4_X1 port map( A1 => n4701, A2 => n4700, A3 => n4699, A4 => 
                           n4698, ZN => n4702);
   U2750 : AOI22_X1 port map( A1 => n4703, A2 => n23, B1 => n4702, B2 => n22, 
                           ZN => n4704);
   U2751 : OAI221_X1 port map( B1 => n5673, B2 => n4706, C1 => n5671, C2 => 
                           n4705, A => n4704, ZN => N271);
   U2752 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n429, B1 => 
                           REGISTERS_23_18_port, B2 => n392, ZN => n4710);
   U2753 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n503, B1 => 
                           REGISTERS_19_18_port, B2 => n466, ZN => n4709);
   U2754 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n577, B1 => 
                           REGISTERS_22_18_port, B2 => n540, ZN => n4708);
   U2755 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n651, B1 => 
                           REGISTERS_18_18_port, B2 => n614, ZN => n4707);
   U2756 : AND4_X1 port map( A1 => n4710, A2 => n4709, A3 => n4708, A4 => n4707
                           , ZN => n4727);
   U2757 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n429, B1 => 
                           REGISTERS_31_18_port, B2 => n392, ZN => n4714);
   U2758 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n503, B1 => 
                           REGISTERS_27_18_port, B2 => n466, ZN => n4713);
   U2759 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n577, B1 => 
                           REGISTERS_30_18_port, B2 => n540, ZN => n4712);
   U2760 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n651, B1 => 
                           REGISTERS_26_18_port, B2 => n614, ZN => n4711);
   U2761 : AND4_X1 port map( A1 => n4714, A2 => n4713, A3 => n4712, A4 => n4711
                           , ZN => n4726);
   U2762 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n429, B1 => 
                           REGISTERS_7_18_port, B2 => n392, ZN => n4718);
   U2763 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n503, B1 => 
                           REGISTERS_3_18_port, B2 => n466, ZN => n4717);
   U2764 : AOI22_X1 port map( A1 => REGISTERS_4_18_port, A2 => n577, B1 => 
                           REGISTERS_6_18_port, B2 => n540, ZN => n4716);
   U2765 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n651, B1 => 
                           REGISTERS_2_18_port, B2 => n614, ZN => n4715);
   U2766 : NAND4_X1 port map( A1 => n4718, A2 => n4717, A3 => n4716, A4 => 
                           n4715, ZN => n4724);
   U2767 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n429, B1 => 
                           REGISTERS_15_18_port, B2 => n392, ZN => n4722);
   U2768 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n503, B1 => 
                           REGISTERS_11_18_port, B2 => n466, ZN => n4721);
   U2769 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n577, B1 => 
                           REGISTERS_14_18_port, B2 => n540, ZN => n4720);
   U2770 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n651, B1 => 
                           REGISTERS_10_18_port, B2 => n614, ZN => n4719);
   U2771 : NAND4_X1 port map( A1 => n4722, A2 => n4721, A3 => n4720, A4 => 
                           n4719, ZN => n4723);
   U2772 : AOI22_X1 port map( A1 => n4724, A2 => n23, B1 => n4723, B2 => n22, 
                           ZN => n4725);
   U2773 : OAI221_X1 port map( B1 => n5673, B2 => n4727, C1 => n5671, C2 => 
                           n4726, A => n4725, ZN => N270);
   U2774 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n429, B1 => 
                           REGISTERS_23_19_port, B2 => n392, ZN => n4731);
   U2775 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n503, B1 => 
                           REGISTERS_19_19_port, B2 => n466, ZN => n4730);
   U2776 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n577, B1 => 
                           REGISTERS_22_19_port, B2 => n540, ZN => n4729);
   U2777 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n651, B1 => 
                           REGISTERS_18_19_port, B2 => n614, ZN => n4728);
   U2778 : AND4_X1 port map( A1 => n4731, A2 => n4730, A3 => n4729, A4 => n4728
                           , ZN => n4748);
   U2779 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n429, B1 => 
                           REGISTERS_31_19_port, B2 => n392, ZN => n4735);
   U2780 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n503, B1 => 
                           REGISTERS_27_19_port, B2 => n466, ZN => n4734);
   U2781 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n577, B1 => 
                           REGISTERS_30_19_port, B2 => n540, ZN => n4733);
   U2782 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n651, B1 => 
                           REGISTERS_26_19_port, B2 => n614, ZN => n4732);
   U2783 : AND4_X1 port map( A1 => n4735, A2 => n4734, A3 => n4733, A4 => n4732
                           , ZN => n4747);
   U2784 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n429, B1 => 
                           REGISTERS_7_19_port, B2 => n392, ZN => n4739);
   U2785 : AOI22_X1 port map( A1 => REGISTERS_1_19_port, A2 => n503, B1 => 
                           REGISTERS_3_19_port, B2 => n466, ZN => n4738);
   U2786 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n577, B1 => 
                           REGISTERS_6_19_port, B2 => n540, ZN => n4737);
   U2787 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n651, B1 => 
                           REGISTERS_2_19_port, B2 => n614, ZN => n4736);
   U2788 : NAND4_X1 port map( A1 => n4739, A2 => n4738, A3 => n4737, A4 => 
                           n4736, ZN => n4745);
   U2789 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n429, B1 => 
                           REGISTERS_15_19_port, B2 => n392, ZN => n4743);
   U2790 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n503, B1 => 
                           REGISTERS_11_19_port, B2 => n466, ZN => n4742);
   U2791 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n577, B1 => 
                           REGISTERS_14_19_port, B2 => n540, ZN => n4741);
   U2792 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n651, B1 => 
                           REGISTERS_10_19_port, B2 => n614, ZN => n4740);
   U2793 : NAND4_X1 port map( A1 => n4743, A2 => n4742, A3 => n4741, A4 => 
                           n4740, ZN => n4744);
   U2794 : AOI22_X1 port map( A1 => n4745, A2 => n23, B1 => n4744, B2 => n22, 
                           ZN => n4746);
   U2795 : OAI221_X1 port map( B1 => n5673, B2 => n4748, C1 => n5671, C2 => 
                           n4747, A => n4746, ZN => N269);
   U2796 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n429, B1 => 
                           REGISTERS_23_20_port, B2 => n392, ZN => n4752);
   U2797 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n503, B1 => 
                           REGISTERS_19_20_port, B2 => n466, ZN => n4751);
   U2798 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n577, B1 => 
                           REGISTERS_22_20_port, B2 => n540, ZN => n4750);
   U2799 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n651, B1 => 
                           REGISTERS_18_20_port, B2 => n614, ZN => n4749);
   U2800 : AND4_X1 port map( A1 => n4752, A2 => n4751, A3 => n4750, A4 => n4749
                           , ZN => n4769);
   U2801 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n429, B1 => 
                           REGISTERS_31_20_port, B2 => n392, ZN => n4756);
   U2802 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n503, B1 => 
                           REGISTERS_27_20_port, B2 => n466, ZN => n4755);
   U2803 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n577, B1 => 
                           REGISTERS_30_20_port, B2 => n540, ZN => n4754);
   U2804 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n651, B1 => 
                           REGISTERS_26_20_port, B2 => n614, ZN => n4753);
   U2805 : AND4_X1 port map( A1 => n4756, A2 => n4755, A3 => n4754, A4 => n4753
                           , ZN => n4768);
   U2806 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n429, B1 => 
                           REGISTERS_7_20_port, B2 => n392, ZN => n4760);
   U2807 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n503, B1 => 
                           REGISTERS_3_20_port, B2 => n466, ZN => n4759);
   U2808 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n577, B1 => 
                           REGISTERS_6_20_port, B2 => n540, ZN => n4758);
   U2809 : AOI22_X1 port map( A1 => REGISTERS_0_20_port, A2 => n651, B1 => 
                           REGISTERS_2_20_port, B2 => n614, ZN => n4757);
   U2810 : NAND4_X1 port map( A1 => n4760, A2 => n4759, A3 => n4758, A4 => 
                           n4757, ZN => n4766);
   U2811 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n429, B1 => 
                           REGISTERS_15_20_port, B2 => n392, ZN => n4764);
   U2812 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n503, B1 => 
                           REGISTERS_11_20_port, B2 => n466, ZN => n4763);
   U2813 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n577, B1 => 
                           REGISTERS_14_20_port, B2 => n540, ZN => n4762);
   U2814 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n651, B1 => 
                           REGISTERS_10_20_port, B2 => n614, ZN => n4761);
   U2815 : NAND4_X1 port map( A1 => n4764, A2 => n4763, A3 => n4762, A4 => 
                           n4761, ZN => n4765);
   U2816 : AOI22_X1 port map( A1 => n4766, A2 => n23, B1 => n4765, B2 => n22, 
                           ZN => n4767);
   U2817 : OAI221_X1 port map( B1 => n5673, B2 => n4769, C1 => n5671, C2 => 
                           n4768, A => n4767, ZN => N268);
   U2818 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n430, B1 => 
                           REGISTERS_23_21_port, B2 => n393, ZN => n4773);
   U2819 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n504, B1 => 
                           REGISTERS_19_21_port, B2 => n467, ZN => n4772);
   U2820 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n578, B1 => 
                           REGISTERS_22_21_port, B2 => n541, ZN => n4771);
   U2821 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n652, B1 => 
                           REGISTERS_18_21_port, B2 => n615, ZN => n4770);
   U2822 : AND4_X1 port map( A1 => n4773, A2 => n4772, A3 => n4771, A4 => n4770
                           , ZN => n4790);
   U2823 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n430, B1 => 
                           REGISTERS_31_21_port, B2 => n393, ZN => n4777);
   U2824 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n504, B1 => 
                           REGISTERS_27_21_port, B2 => n467, ZN => n4776);
   U2825 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n578, B1 => 
                           REGISTERS_30_21_port, B2 => n541, ZN => n4775);
   U2826 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n652, B1 => 
                           REGISTERS_26_21_port, B2 => n615, ZN => n4774);
   U2827 : AND4_X1 port map( A1 => n4777, A2 => n4776, A3 => n4775, A4 => n4774
                           , ZN => n4789);
   U2828 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n430, B1 => 
                           REGISTERS_7_21_port, B2 => n393, ZN => n4781);
   U2829 : AOI22_X1 port map( A1 => REGISTERS_1_21_port, A2 => n504, B1 => 
                           REGISTERS_3_21_port, B2 => n467, ZN => n4780);
   U2830 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n578, B1 => 
                           REGISTERS_6_21_port, B2 => n541, ZN => n4779);
   U2831 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n652, B1 => 
                           REGISTERS_2_21_port, B2 => n615, ZN => n4778);
   U2832 : NAND4_X1 port map( A1 => n4781, A2 => n4780, A3 => n4779, A4 => 
                           n4778, ZN => n4787);
   U2833 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n430, B1 => 
                           REGISTERS_15_21_port, B2 => n393, ZN => n4785);
   U2834 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n504, B1 => 
                           REGISTERS_11_21_port, B2 => n467, ZN => n4784);
   U2835 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n578, B1 => 
                           REGISTERS_14_21_port, B2 => n541, ZN => n4783);
   U2836 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n652, B1 => 
                           REGISTERS_10_21_port, B2 => n615, ZN => n4782);
   U2837 : NAND4_X1 port map( A1 => n4785, A2 => n4784, A3 => n4783, A4 => 
                           n4782, ZN => n4786);
   U2838 : AOI22_X1 port map( A1 => n4787, A2 => n23, B1 => n4786, B2 => n22, 
                           ZN => n4788);
   U2839 : OAI221_X1 port map( B1 => n5673, B2 => n4790, C1 => n5671, C2 => 
                           n4789, A => n4788, ZN => N267);
   U2840 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n430, B1 => 
                           REGISTERS_23_22_port, B2 => n393, ZN => n4794);
   U2841 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n504, B1 => 
                           REGISTERS_19_22_port, B2 => n467, ZN => n4793);
   U2842 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n578, B1 => 
                           REGISTERS_22_22_port, B2 => n541, ZN => n4792);
   U2843 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n652, B1 => 
                           REGISTERS_18_22_port, B2 => n615, ZN => n4791);
   U2844 : AND4_X1 port map( A1 => n4794, A2 => n4793, A3 => n4792, A4 => n4791
                           , ZN => n4811);
   U2845 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n430, B1 => 
                           REGISTERS_31_22_port, B2 => n393, ZN => n4798);
   U2846 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n504, B1 => 
                           REGISTERS_27_22_port, B2 => n467, ZN => n4797);
   U2847 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n578, B1 => 
                           REGISTERS_30_22_port, B2 => n541, ZN => n4796);
   U2848 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n652, B1 => 
                           REGISTERS_26_22_port, B2 => n615, ZN => n4795);
   U2849 : AND4_X1 port map( A1 => n4798, A2 => n4797, A3 => n4796, A4 => n4795
                           , ZN => n4810);
   U2850 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n430, B1 => 
                           REGISTERS_7_22_port, B2 => n393, ZN => n4802);
   U2851 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n504, B1 => 
                           REGISTERS_3_22_port, B2 => n467, ZN => n4801);
   U2852 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n578, B1 => 
                           REGISTERS_6_22_port, B2 => n541, ZN => n4800);
   U2853 : AOI22_X1 port map( A1 => REGISTERS_0_22_port, A2 => n652, B1 => 
                           REGISTERS_2_22_port, B2 => n615, ZN => n4799);
   U2854 : NAND4_X1 port map( A1 => n4802, A2 => n4801, A3 => n4800, A4 => 
                           n4799, ZN => n4808);
   U2855 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n430, B1 => 
                           REGISTERS_15_22_port, B2 => n393, ZN => n4806);
   U2856 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n504, B1 => 
                           REGISTERS_11_22_port, B2 => n467, ZN => n4805);
   U2857 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n578, B1 => 
                           REGISTERS_14_22_port, B2 => n541, ZN => n4804);
   U2858 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n652, B1 => 
                           REGISTERS_10_22_port, B2 => n615, ZN => n4803);
   U2859 : NAND4_X1 port map( A1 => n4806, A2 => n4805, A3 => n4804, A4 => 
                           n4803, ZN => n4807);
   U2860 : AOI22_X1 port map( A1 => n4808, A2 => n23, B1 => n4807, B2 => n22, 
                           ZN => n4809);
   U2861 : OAI221_X1 port map( B1 => n5673, B2 => n4811, C1 => n5671, C2 => 
                           n4810, A => n4809, ZN => N266);
   U2862 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n430, B1 => 
                           REGISTERS_23_23_port, B2 => n393, ZN => n4815);
   U2863 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n504, B1 => 
                           REGISTERS_19_23_port, B2 => n467, ZN => n4814);
   U2864 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n578, B1 => 
                           REGISTERS_22_23_port, B2 => n541, ZN => n4813);
   U2865 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n652, B1 => 
                           REGISTERS_18_23_port, B2 => n615, ZN => n4812);
   U2866 : AND4_X1 port map( A1 => n4815, A2 => n4814, A3 => n4813, A4 => n4812
                           , ZN => n4832);
   U2867 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n430, B1 => 
                           REGISTERS_31_23_port, B2 => n393, ZN => n4819);
   U2868 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n504, B1 => 
                           REGISTERS_27_23_port, B2 => n467, ZN => n4818);
   U2869 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n578, B1 => 
                           REGISTERS_30_23_port, B2 => n541, ZN => n4817);
   U2870 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n652, B1 => 
                           REGISTERS_26_23_port, B2 => n615, ZN => n4816);
   U2871 : AND4_X1 port map( A1 => n4819, A2 => n4818, A3 => n4817, A4 => n4816
                           , ZN => n4831);
   U2872 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n430, B1 => 
                           REGISTERS_7_23_port, B2 => n393, ZN => n4823);
   U2873 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n504, B1 => 
                           REGISTERS_3_23_port, B2 => n467, ZN => n4822);
   U2874 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n578, B1 => 
                           REGISTERS_6_23_port, B2 => n541, ZN => n4821);
   U2875 : AOI22_X1 port map( A1 => REGISTERS_0_23_port, A2 => n652, B1 => 
                           REGISTERS_2_23_port, B2 => n615, ZN => n4820);
   U2876 : NAND4_X1 port map( A1 => n4823, A2 => n4822, A3 => n4821, A4 => 
                           n4820, ZN => n4829);
   U2877 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n430, B1 => 
                           REGISTERS_15_23_port, B2 => n393, ZN => n4827);
   U2878 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n504, B1 => 
                           REGISTERS_11_23_port, B2 => n467, ZN => n4826);
   U2879 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n578, B1 => 
                           REGISTERS_14_23_port, B2 => n541, ZN => n4825);
   U2880 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n652, B1 => 
                           REGISTERS_10_23_port, B2 => n615, ZN => n4824);
   U2881 : NAND4_X1 port map( A1 => n4827, A2 => n4826, A3 => n4825, A4 => 
                           n4824, ZN => n4828);
   U2882 : AOI22_X1 port map( A1 => n4829, A2 => n23, B1 => n4828, B2 => n22, 
                           ZN => n4830);
   U2883 : OAI221_X1 port map( B1 => n5673, B2 => n4832, C1 => n5671, C2 => 
                           n4831, A => n4830, ZN => N265);
   U2884 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n431, B1 => 
                           REGISTERS_23_24_port, B2 => n394, ZN => n4836);
   U2885 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n505, B1 => 
                           REGISTERS_19_24_port, B2 => n468, ZN => n4835);
   U2886 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n579, B1 => 
                           REGISTERS_22_24_port, B2 => n542, ZN => n4834);
   U2887 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n653, B1 => 
                           REGISTERS_18_24_port, B2 => n616, ZN => n4833);
   U2888 : AND4_X1 port map( A1 => n4836, A2 => n4835, A3 => n4834, A4 => n4833
                           , ZN => n4853);
   U2889 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n431, B1 => 
                           REGISTERS_31_24_port, B2 => n394, ZN => n4840);
   U2890 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n505, B1 => 
                           REGISTERS_27_24_port, B2 => n468, ZN => n4839);
   U2891 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n579, B1 => 
                           REGISTERS_30_24_port, B2 => n542, ZN => n4838);
   U2892 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n653, B1 => 
                           REGISTERS_26_24_port, B2 => n616, ZN => n4837);
   U2893 : AND4_X1 port map( A1 => n4840, A2 => n4839, A3 => n4838, A4 => n4837
                           , ZN => n4852);
   U2894 : AOI22_X1 port map( A1 => REGISTERS_5_24_port, A2 => n431, B1 => 
                           REGISTERS_7_24_port, B2 => n394, ZN => n4844);
   U2895 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n505, B1 => 
                           REGISTERS_3_24_port, B2 => n468, ZN => n4843);
   U2896 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n579, B1 => 
                           REGISTERS_6_24_port, B2 => n542, ZN => n4842);
   U2897 : AOI22_X1 port map( A1 => REGISTERS_0_24_port, A2 => n653, B1 => 
                           REGISTERS_2_24_port, B2 => n616, ZN => n4841);
   U2898 : NAND4_X1 port map( A1 => n4844, A2 => n4843, A3 => n4842, A4 => 
                           n4841, ZN => n4850);
   U2899 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n431, B1 => 
                           REGISTERS_15_24_port, B2 => n394, ZN => n4848);
   U2900 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n505, B1 => 
                           REGISTERS_11_24_port, B2 => n468, ZN => n4847);
   U2901 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n579, B1 => 
                           REGISTERS_14_24_port, B2 => n542, ZN => n4846);
   U2902 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n653, B1 => 
                           REGISTERS_10_24_port, B2 => n616, ZN => n4845);
   U2903 : NAND4_X1 port map( A1 => n4848, A2 => n4847, A3 => n4846, A4 => 
                           n4845, ZN => n4849);
   U2904 : AOI22_X1 port map( A1 => n4850, A2 => n23, B1 => n4849, B2 => n22, 
                           ZN => n4851);
   U2905 : OAI221_X1 port map( B1 => n5673, B2 => n4853, C1 => n5671, C2 => 
                           n4852, A => n4851, ZN => N264);
   U2906 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n431, B1 => 
                           REGISTERS_23_25_port, B2 => n394, ZN => n4857);
   U2907 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n505, B1 => 
                           REGISTERS_19_25_port, B2 => n468, ZN => n4856);
   U2908 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n579, B1 => 
                           REGISTERS_22_25_port, B2 => n542, ZN => n4855);
   U2909 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n653, B1 => 
                           REGISTERS_18_25_port, B2 => n616, ZN => n4854);
   U2910 : AND4_X1 port map( A1 => n4857, A2 => n4856, A3 => n4855, A4 => n4854
                           , ZN => n4874);
   U2911 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n431, B1 => 
                           REGISTERS_31_25_port, B2 => n394, ZN => n4861);
   U2912 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n505, B1 => 
                           REGISTERS_27_25_port, B2 => n468, ZN => n4860);
   U2913 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n579, B1 => 
                           REGISTERS_30_25_port, B2 => n542, ZN => n4859);
   U2914 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n653, B1 => 
                           REGISTERS_26_25_port, B2 => n616, ZN => n4858);
   U2915 : AND4_X1 port map( A1 => n4861, A2 => n4860, A3 => n4859, A4 => n4858
                           , ZN => n4873);
   U2916 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n431, B1 => 
                           REGISTERS_7_25_port, B2 => n394, ZN => n4865);
   U2917 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n505, B1 => 
                           REGISTERS_3_25_port, B2 => n468, ZN => n4864);
   U2918 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n579, B1 => 
                           REGISTERS_6_25_port, B2 => n542, ZN => n4863);
   U2919 : AOI22_X1 port map( A1 => REGISTERS_0_25_port, A2 => n653, B1 => 
                           REGISTERS_2_25_port, B2 => n616, ZN => n4862);
   U2920 : NAND4_X1 port map( A1 => n4865, A2 => n4864, A3 => n4863, A4 => 
                           n4862, ZN => n4871);
   U2921 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n431, B1 => 
                           REGISTERS_15_25_port, B2 => n394, ZN => n4869);
   U2922 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n505, B1 => 
                           REGISTERS_11_25_port, B2 => n468, ZN => n4868);
   U2923 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n579, B1 => 
                           REGISTERS_14_25_port, B2 => n542, ZN => n4867);
   U2924 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n653, B1 => 
                           REGISTERS_10_25_port, B2 => n616, ZN => n4866);
   U2925 : NAND4_X1 port map( A1 => n4869, A2 => n4868, A3 => n4867, A4 => 
                           n4866, ZN => n4870);
   U2926 : AOI22_X1 port map( A1 => n4871, A2 => n23, B1 => n4870, B2 => n22, 
                           ZN => n4872);
   U2927 : OAI221_X1 port map( B1 => n5673, B2 => n4874, C1 => n5671, C2 => 
                           n4873, A => n4872, ZN => N263);
   U2928 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n431, B1 => 
                           REGISTERS_23_26_port, B2 => n394, ZN => n4878);
   U2929 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n505, B1 => 
                           REGISTERS_19_26_port, B2 => n468, ZN => n4877);
   U2930 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n579, B1 => 
                           REGISTERS_22_26_port, B2 => n542, ZN => n4876);
   U2931 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n653, B1 => 
                           REGISTERS_18_26_port, B2 => n616, ZN => n4875);
   U2932 : AND4_X1 port map( A1 => n4878, A2 => n4877, A3 => n4876, A4 => n4875
                           , ZN => n4895);
   U2933 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n431, B1 => 
                           REGISTERS_31_26_port, B2 => n394, ZN => n4882);
   U2934 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n505, B1 => 
                           REGISTERS_27_26_port, B2 => n468, ZN => n4881);
   U2935 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n579, B1 => 
                           REGISTERS_30_26_port, B2 => n542, ZN => n4880);
   U2936 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n653, B1 => 
                           REGISTERS_26_26_port, B2 => n616, ZN => n4879);
   U2937 : AND4_X1 port map( A1 => n4882, A2 => n4881, A3 => n4880, A4 => n4879
                           , ZN => n4894);
   U2938 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n431, B1 => 
                           REGISTERS_7_26_port, B2 => n394, ZN => n4886);
   U2939 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n505, B1 => 
                           REGISTERS_3_26_port, B2 => n468, ZN => n4885);
   U2940 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n579, B1 => 
                           REGISTERS_6_26_port, B2 => n542, ZN => n4884);
   U2941 : AOI22_X1 port map( A1 => REGISTERS_0_26_port, A2 => n653, B1 => 
                           REGISTERS_2_26_port, B2 => n616, ZN => n4883);
   U2942 : NAND4_X1 port map( A1 => n4886, A2 => n4885, A3 => n4884, A4 => 
                           n4883, ZN => n4892);
   U2943 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n431, B1 => 
                           REGISTERS_15_26_port, B2 => n394, ZN => n4890);
   U2944 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n505, B1 => 
                           REGISTERS_11_26_port, B2 => n468, ZN => n4889);
   U2945 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n579, B1 => 
                           REGISTERS_14_26_port, B2 => n542, ZN => n4888);
   U2946 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n653, B1 => 
                           REGISTERS_10_26_port, B2 => n616, ZN => n4887);
   U2947 : NAND4_X1 port map( A1 => n4890, A2 => n4889, A3 => n4888, A4 => 
                           n4887, ZN => n4891);
   U2948 : AOI22_X1 port map( A1 => n4892, A2 => n23, B1 => n4891, B2 => n22, 
                           ZN => n4893);
   U2949 : OAI221_X1 port map( B1 => n5673, B2 => n4895, C1 => n5671, C2 => 
                           n4894, A => n4893, ZN => N262);
   U2950 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n432, B1 => 
                           REGISTERS_23_27_port, B2 => n395, ZN => n4899);
   U2951 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n506, B1 => 
                           REGISTERS_19_27_port, B2 => n469, ZN => n4898);
   U2952 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n580, B1 => 
                           REGISTERS_22_27_port, B2 => n543, ZN => n4897);
   U2953 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n654, B1 => 
                           REGISTERS_18_27_port, B2 => n617, ZN => n4896);
   U2954 : AND4_X1 port map( A1 => n4899, A2 => n4898, A3 => n4897, A4 => n4896
                           , ZN => n4916);
   U2955 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n432, B1 => 
                           REGISTERS_31_27_port, B2 => n395, ZN => n4903);
   U2956 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n506, B1 => 
                           REGISTERS_27_27_port, B2 => n469, ZN => n4902);
   U2957 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n580, B1 => 
                           REGISTERS_30_27_port, B2 => n543, ZN => n4901);
   U2958 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n654, B1 => 
                           REGISTERS_26_27_port, B2 => n617, ZN => n4900);
   U2959 : AND4_X1 port map( A1 => n4903, A2 => n4902, A3 => n4901, A4 => n4900
                           , ZN => n4915);
   U2960 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n432, B1 => 
                           REGISTERS_7_27_port, B2 => n395, ZN => n4907);
   U2961 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n506, B1 => 
                           REGISTERS_3_27_port, B2 => n469, ZN => n4906);
   U2962 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n580, B1 => 
                           REGISTERS_6_27_port, B2 => n543, ZN => n4905);
   U2963 : AOI22_X1 port map( A1 => REGISTERS_0_27_port, A2 => n654, B1 => 
                           REGISTERS_2_27_port, B2 => n617, ZN => n4904);
   U2964 : NAND4_X1 port map( A1 => n4907, A2 => n4906, A3 => n4905, A4 => 
                           n4904, ZN => n4913);
   U2965 : AOI22_X1 port map( A1 => REGISTERS_13_27_port, A2 => n432, B1 => 
                           REGISTERS_15_27_port, B2 => n395, ZN => n4911);
   U2966 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n506, B1 => 
                           REGISTERS_11_27_port, B2 => n469, ZN => n4910);
   U2967 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n580, B1 => 
                           REGISTERS_14_27_port, B2 => n543, ZN => n4909);
   U2968 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n654, B1 => 
                           REGISTERS_10_27_port, B2 => n617, ZN => n4908);
   U2969 : NAND4_X1 port map( A1 => n4911, A2 => n4910, A3 => n4909, A4 => 
                           n4908, ZN => n4912);
   U2970 : AOI22_X1 port map( A1 => n4913, A2 => n23, B1 => n4912, B2 => n22, 
                           ZN => n4914);
   U2971 : OAI221_X1 port map( B1 => n5673, B2 => n4916, C1 => n5671, C2 => 
                           n4915, A => n4914, ZN => N261);
   U2972 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n432, B1 => 
                           REGISTERS_23_28_port, B2 => n395, ZN => n4920);
   U2973 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n506, B1 => 
                           REGISTERS_19_28_port, B2 => n469, ZN => n4919);
   U2974 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n580, B1 => 
                           REGISTERS_22_28_port, B2 => n543, ZN => n4918);
   U2975 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n654, B1 => 
                           REGISTERS_18_28_port, B2 => n617, ZN => n4917);
   U2976 : AND4_X1 port map( A1 => n4920, A2 => n4919, A3 => n4918, A4 => n4917
                           , ZN => n4937);
   U2977 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n432, B1 => 
                           REGISTERS_31_28_port, B2 => n395, ZN => n4924);
   U2978 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n506, B1 => 
                           REGISTERS_27_28_port, B2 => n469, ZN => n4923);
   U2979 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n580, B1 => 
                           REGISTERS_30_28_port, B2 => n543, ZN => n4922);
   U2980 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n654, B1 => 
                           REGISTERS_26_28_port, B2 => n617, ZN => n4921);
   U2981 : AND4_X1 port map( A1 => n4924, A2 => n4923, A3 => n4922, A4 => n4921
                           , ZN => n4936);
   U2982 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n432, B1 => 
                           REGISTERS_7_28_port, B2 => n395, ZN => n4928);
   U2983 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n506, B1 => 
                           REGISTERS_3_28_port, B2 => n469, ZN => n4927);
   U2984 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n580, B1 => 
                           REGISTERS_6_28_port, B2 => n543, ZN => n4926);
   U2985 : AOI22_X1 port map( A1 => REGISTERS_0_28_port, A2 => n654, B1 => 
                           REGISTERS_2_28_port, B2 => n617, ZN => n4925);
   U2986 : NAND4_X1 port map( A1 => n4928, A2 => n4927, A3 => n4926, A4 => 
                           n4925, ZN => n4934);
   U2987 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n432, B1 => 
                           REGISTERS_15_28_port, B2 => n395, ZN => n4932);
   U2988 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n506, B1 => 
                           REGISTERS_11_28_port, B2 => n469, ZN => n4931);
   U2989 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n580, B1 => 
                           REGISTERS_14_28_port, B2 => n543, ZN => n4930);
   U2990 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n654, B1 => 
                           REGISTERS_10_28_port, B2 => n617, ZN => n4929);
   U2991 : NAND4_X1 port map( A1 => n4932, A2 => n4931, A3 => n4930, A4 => 
                           n4929, ZN => n4933);
   U2992 : AOI22_X1 port map( A1 => n4934, A2 => n23, B1 => n4933, B2 => n22, 
                           ZN => n4935);
   U2993 : OAI221_X1 port map( B1 => n5673, B2 => n4937, C1 => n5671, C2 => 
                           n4936, A => n4935, ZN => N260);
   U2994 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n432, B1 => 
                           REGISTERS_23_29_port, B2 => n395, ZN => n4941);
   U2995 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n506, B1 => 
                           REGISTERS_19_29_port, B2 => n469, ZN => n4940);
   U2996 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n580, B1 => 
                           REGISTERS_22_29_port, B2 => n543, ZN => n4939);
   U2997 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n654, B1 => 
                           REGISTERS_18_29_port, B2 => n617, ZN => n4938);
   U2998 : AND4_X1 port map( A1 => n4941, A2 => n4940, A3 => n4939, A4 => n4938
                           , ZN => n4958);
   U2999 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n432, B1 => 
                           REGISTERS_31_29_port, B2 => n395, ZN => n4945);
   U3000 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n506, B1 => 
                           REGISTERS_27_29_port, B2 => n469, ZN => n4944);
   U3001 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n580, B1 => 
                           REGISTERS_30_29_port, B2 => n543, ZN => n4943);
   U3002 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n654, B1 => 
                           REGISTERS_26_29_port, B2 => n617, ZN => n4942);
   U3003 : AND4_X1 port map( A1 => n4945, A2 => n4944, A3 => n4943, A4 => n4942
                           , ZN => n4957);
   U3004 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n432, B1 => 
                           REGISTERS_7_29_port, B2 => n395, ZN => n4949);
   U3005 : AOI22_X1 port map( A1 => REGISTERS_1_29_port, A2 => n506, B1 => 
                           REGISTERS_3_29_port, B2 => n469, ZN => n4948);
   U3006 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n580, B1 => 
                           REGISTERS_6_29_port, B2 => n543, ZN => n4947);
   U3007 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n654, B1 => 
                           REGISTERS_2_29_port, B2 => n617, ZN => n4946);
   U3008 : NAND4_X1 port map( A1 => n4949, A2 => n4948, A3 => n4947, A4 => 
                           n4946, ZN => n4955);
   U3009 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n432, B1 => 
                           REGISTERS_15_29_port, B2 => n395, ZN => n4953);
   U3010 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n506, B1 => 
                           REGISTERS_11_29_port, B2 => n469, ZN => n4952);
   U3011 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n580, B1 => 
                           REGISTERS_14_29_port, B2 => n543, ZN => n4951);
   U3012 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n654, B1 => 
                           REGISTERS_10_29_port, B2 => n617, ZN => n4950);
   U3013 : NAND4_X1 port map( A1 => n4953, A2 => n4952, A3 => n4951, A4 => 
                           n4950, ZN => n4954);
   U3014 : AOI22_X1 port map( A1 => n4955, A2 => n23, B1 => n4954, B2 => n22, 
                           ZN => n4956);
   U3015 : OAI221_X1 port map( B1 => n5673, B2 => n4958, C1 => n5671, C2 => 
                           n4957, A => n4956, ZN => N259);
   U3016 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n433, B1 => 
                           REGISTERS_23_30_port, B2 => n396, ZN => n4962);
   U3017 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n507, B1 => 
                           REGISTERS_19_30_port, B2 => n470, ZN => n4961);
   U3018 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n581, B1 => 
                           REGISTERS_22_30_port, B2 => n544, ZN => n4960);
   U3019 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n655, B1 => 
                           REGISTERS_18_30_port, B2 => n618, ZN => n4959);
   U3020 : AND4_X1 port map( A1 => n4962, A2 => n4961, A3 => n4960, A4 => n4959
                           , ZN => n4979);
   U3021 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n433, B1 => 
                           REGISTERS_31_30_port, B2 => n396, ZN => n4966);
   U3022 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n507, B1 => 
                           REGISTERS_27_30_port, B2 => n470, ZN => n4965);
   U3023 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n581, B1 => 
                           REGISTERS_30_30_port, B2 => n544, ZN => n4964);
   U3024 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n655, B1 => 
                           REGISTERS_26_30_port, B2 => n618, ZN => n4963);
   U3025 : AND4_X1 port map( A1 => n4966, A2 => n4965, A3 => n4964, A4 => n4963
                           , ZN => n4978);
   U3026 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n433, B1 => 
                           REGISTERS_7_30_port, B2 => n396, ZN => n4970);
   U3027 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n507, B1 => 
                           REGISTERS_3_30_port, B2 => n470, ZN => n4969);
   U3028 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n581, B1 => 
                           REGISTERS_6_30_port, B2 => n544, ZN => n4968);
   U3029 : AOI22_X1 port map( A1 => REGISTERS_0_30_port, A2 => n655, B1 => 
                           REGISTERS_2_30_port, B2 => n618, ZN => n4967);
   U3030 : NAND4_X1 port map( A1 => n4970, A2 => n4969, A3 => n4968, A4 => 
                           n4967, ZN => n4976);
   U3031 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n433, B1 => 
                           REGISTERS_15_30_port, B2 => n396, ZN => n4974);
   U3032 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n507, B1 => 
                           REGISTERS_11_30_port, B2 => n470, ZN => n4973);
   U3033 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n581, B1 => 
                           REGISTERS_14_30_port, B2 => n544, ZN => n4972);
   U3034 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n655, B1 => 
                           REGISTERS_10_30_port, B2 => n618, ZN => n4971);
   U3035 : NAND4_X1 port map( A1 => n4974, A2 => n4973, A3 => n4972, A4 => 
                           n4971, ZN => n4975);
   U3036 : AOI22_X1 port map( A1 => n4976, A2 => n23, B1 => n4975, B2 => n22, 
                           ZN => n4977);
   U3037 : OAI221_X1 port map( B1 => n5673, B2 => n4979, C1 => n5671, C2 => 
                           n4978, A => n4977, ZN => N258);
   U3038 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n433, B1 => 
                           REGISTERS_23_31_port, B2 => n396, ZN => n4983);
   U3039 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n507, B1 => 
                           REGISTERS_19_31_port, B2 => n470, ZN => n4982);
   U3040 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n581, B1 => 
                           REGISTERS_22_31_port, B2 => n544, ZN => n4981);
   U3041 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n655, B1 => 
                           REGISTERS_18_31_port, B2 => n618, ZN => n4980);
   U3042 : AND4_X1 port map( A1 => n4983, A2 => n4982, A3 => n4981, A4 => n4980
                           , ZN => n5000);
   U3043 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n433, B1 => 
                           REGISTERS_31_31_port, B2 => n396, ZN => n4987);
   U3044 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n507, B1 => 
                           REGISTERS_27_31_port, B2 => n470, ZN => n4986);
   U3045 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n581, B1 => 
                           REGISTERS_30_31_port, B2 => n544, ZN => n4985);
   U3046 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n655, B1 => 
                           REGISTERS_26_31_port, B2 => n618, ZN => n4984);
   U3047 : AND4_X1 port map( A1 => n4987, A2 => n4986, A3 => n4985, A4 => n4984
                           , ZN => n4999);
   U3048 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n433, B1 => 
                           REGISTERS_7_31_port, B2 => n396, ZN => n4991);
   U3049 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n507, B1 => 
                           REGISTERS_3_31_port, B2 => n470, ZN => n4990);
   U3050 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n581, B1 => 
                           REGISTERS_6_31_port, B2 => n544, ZN => n4989);
   U3051 : AOI22_X1 port map( A1 => REGISTERS_0_31_port, A2 => n655, B1 => 
                           REGISTERS_2_31_port, B2 => n618, ZN => n4988);
   U3052 : NAND4_X1 port map( A1 => n4991, A2 => n4990, A3 => n4989, A4 => 
                           n4988, ZN => n4997);
   U3053 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n433, B1 => 
                           REGISTERS_15_31_port, B2 => n396, ZN => n4995);
   U3054 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n507, B1 => 
                           REGISTERS_11_31_port, B2 => n470, ZN => n4994);
   U3055 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n581, B1 => 
                           REGISTERS_14_31_port, B2 => n544, ZN => n4993);
   U3056 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n655, B1 => 
                           REGISTERS_10_31_port, B2 => n618, ZN => n4992);
   U3057 : NAND4_X1 port map( A1 => n4995, A2 => n4994, A3 => n4993, A4 => 
                           n4992, ZN => n4996);
   U3058 : AOI22_X1 port map( A1 => n4997, A2 => n23, B1 => n4996, B2 => n22, 
                           ZN => n4998);
   U3059 : OAI221_X1 port map( B1 => n5673, B2 => n5000, C1 => n5671, C2 => 
                           n4999, A => n4998, ZN => N257);
   U3060 : AOI22_X1 port map( A1 => REGISTERS_21_32_port, A2 => n433, B1 => 
                           REGISTERS_23_32_port, B2 => n396, ZN => n5004);
   U3061 : AOI22_X1 port map( A1 => REGISTERS_17_32_port, A2 => n507, B1 => 
                           REGISTERS_19_32_port, B2 => n470, ZN => n5003);
   U3062 : AOI22_X1 port map( A1 => REGISTERS_20_32_port, A2 => n581, B1 => 
                           REGISTERS_22_32_port, B2 => n544, ZN => n5002);
   U3063 : AOI22_X1 port map( A1 => REGISTERS_16_32_port, A2 => n655, B1 => 
                           REGISTERS_18_32_port, B2 => n618, ZN => n5001);
   U3064 : AND4_X1 port map( A1 => n5004, A2 => n5003, A3 => n5002, A4 => n5001
                           , ZN => n5021);
   U3065 : AOI22_X1 port map( A1 => REGISTERS_29_32_port, A2 => n433, B1 => 
                           REGISTERS_31_32_port, B2 => n396, ZN => n5008);
   U3066 : AOI22_X1 port map( A1 => REGISTERS_25_32_port, A2 => n507, B1 => 
                           REGISTERS_27_32_port, B2 => n470, ZN => n5007);
   U3067 : AOI22_X1 port map( A1 => REGISTERS_28_32_port, A2 => n581, B1 => 
                           REGISTERS_30_32_port, B2 => n544, ZN => n5006);
   U3068 : AOI22_X1 port map( A1 => REGISTERS_24_32_port, A2 => n655, B1 => 
                           REGISTERS_26_32_port, B2 => n618, ZN => n5005);
   U3069 : AND4_X1 port map( A1 => n5008, A2 => n5007, A3 => n5006, A4 => n5005
                           , ZN => n5020);
   U3070 : AOI22_X1 port map( A1 => REGISTERS_5_32_port, A2 => n433, B1 => 
                           REGISTERS_7_32_port, B2 => n396, ZN => n5012);
   U3071 : AOI22_X1 port map( A1 => REGISTERS_1_32_port, A2 => n507, B1 => 
                           REGISTERS_3_32_port, B2 => n470, ZN => n5011);
   U3072 : AOI22_X1 port map( A1 => REGISTERS_4_32_port, A2 => n581, B1 => 
                           REGISTERS_6_32_port, B2 => n544, ZN => n5010);
   U3073 : AOI22_X1 port map( A1 => REGISTERS_0_32_port, A2 => n655, B1 => 
                           REGISTERS_2_32_port, B2 => n618, ZN => n5009);
   U3074 : NAND4_X1 port map( A1 => n5012, A2 => n5011, A3 => n5010, A4 => 
                           n5009, ZN => n5018);
   U3075 : AOI22_X1 port map( A1 => REGISTERS_13_32_port, A2 => n433, B1 => 
                           REGISTERS_15_32_port, B2 => n396, ZN => n5016);
   U3076 : AOI22_X1 port map( A1 => REGISTERS_9_32_port, A2 => n507, B1 => 
                           REGISTERS_11_32_port, B2 => n470, ZN => n5015);
   U3077 : AOI22_X1 port map( A1 => REGISTERS_12_32_port, A2 => n581, B1 => 
                           REGISTERS_14_32_port, B2 => n544, ZN => n5014);
   U3078 : AOI22_X1 port map( A1 => REGISTERS_8_32_port, A2 => n655, B1 => 
                           REGISTERS_10_32_port, B2 => n618, ZN => n5013);
   U3079 : NAND4_X1 port map( A1 => n5016, A2 => n5015, A3 => n5014, A4 => 
                           n5013, ZN => n5017);
   U3080 : AOI22_X1 port map( A1 => n5018, A2 => n23, B1 => n5017, B2 => n22, 
                           ZN => n5019);
   U3081 : OAI221_X1 port map( B1 => n5673, B2 => n5021, C1 => n5671, C2 => 
                           n5020, A => n5019, ZN => N256);
   U3082 : AOI22_X1 port map( A1 => REGISTERS_21_33_port, A2 => n434, B1 => 
                           REGISTERS_23_33_port, B2 => n397, ZN => n5025);
   U3083 : AOI22_X1 port map( A1 => REGISTERS_17_33_port, A2 => n508, B1 => 
                           REGISTERS_19_33_port, B2 => n471, ZN => n5024);
   U3084 : AOI22_X1 port map( A1 => REGISTERS_20_33_port, A2 => n582, B1 => 
                           REGISTERS_22_33_port, B2 => n545, ZN => n5023);
   U3085 : AOI22_X1 port map( A1 => REGISTERS_16_33_port, A2 => n656, B1 => 
                           REGISTERS_18_33_port, B2 => n619, ZN => n5022);
   U3086 : AND4_X1 port map( A1 => n5025, A2 => n5024, A3 => n5023, A4 => n5022
                           , ZN => n5042);
   U3087 : AOI22_X1 port map( A1 => REGISTERS_29_33_port, A2 => n434, B1 => 
                           REGISTERS_31_33_port, B2 => n397, ZN => n5029);
   U3088 : AOI22_X1 port map( A1 => REGISTERS_25_33_port, A2 => n508, B1 => 
                           REGISTERS_27_33_port, B2 => n471, ZN => n5028);
   U3089 : AOI22_X1 port map( A1 => REGISTERS_28_33_port, A2 => n582, B1 => 
                           REGISTERS_30_33_port, B2 => n545, ZN => n5027);
   U3090 : AOI22_X1 port map( A1 => REGISTERS_24_33_port, A2 => n656, B1 => 
                           REGISTERS_26_33_port, B2 => n619, ZN => n5026);
   U3091 : AND4_X1 port map( A1 => n5029, A2 => n5028, A3 => n5027, A4 => n5026
                           , ZN => n5041);
   U3092 : AOI22_X1 port map( A1 => REGISTERS_5_33_port, A2 => n434, B1 => 
                           REGISTERS_7_33_port, B2 => n397, ZN => n5033);
   U3093 : AOI22_X1 port map( A1 => REGISTERS_1_33_port, A2 => n508, B1 => 
                           REGISTERS_3_33_port, B2 => n471, ZN => n5032);
   U3094 : AOI22_X1 port map( A1 => REGISTERS_4_33_port, A2 => n582, B1 => 
                           REGISTERS_6_33_port, B2 => n545, ZN => n5031);
   U3095 : AOI22_X1 port map( A1 => REGISTERS_0_33_port, A2 => n656, B1 => 
                           REGISTERS_2_33_port, B2 => n619, ZN => n5030);
   U3096 : NAND4_X1 port map( A1 => n5033, A2 => n5032, A3 => n5031, A4 => 
                           n5030, ZN => n5039);
   U3097 : AOI22_X1 port map( A1 => REGISTERS_13_33_port, A2 => n434, B1 => 
                           REGISTERS_15_33_port, B2 => n397, ZN => n5037);
   U3098 : AOI22_X1 port map( A1 => REGISTERS_9_33_port, A2 => n508, B1 => 
                           REGISTERS_11_33_port, B2 => n471, ZN => n5036);
   U3099 : AOI22_X1 port map( A1 => REGISTERS_12_33_port, A2 => n582, B1 => 
                           REGISTERS_14_33_port, B2 => n545, ZN => n5035);
   U3100 : AOI22_X1 port map( A1 => REGISTERS_8_33_port, A2 => n656, B1 => 
                           REGISTERS_10_33_port, B2 => n619, ZN => n5034);
   U3101 : NAND4_X1 port map( A1 => n5037, A2 => n5036, A3 => n5035, A4 => 
                           n5034, ZN => n5038);
   U3102 : AOI22_X1 port map( A1 => n5039, A2 => n23, B1 => n5038, B2 => n22, 
                           ZN => n5040);
   U3103 : OAI221_X1 port map( B1 => n5673, B2 => n5042, C1 => n5671, C2 => 
                           n5041, A => n5040, ZN => N255);
   U3104 : AOI22_X1 port map( A1 => REGISTERS_21_34_port, A2 => n434, B1 => 
                           REGISTERS_23_34_port, B2 => n397, ZN => n5046);
   U3105 : AOI22_X1 port map( A1 => REGISTERS_17_34_port, A2 => n508, B1 => 
                           REGISTERS_19_34_port, B2 => n471, ZN => n5045);
   U3106 : AOI22_X1 port map( A1 => REGISTERS_20_34_port, A2 => n582, B1 => 
                           REGISTERS_22_34_port, B2 => n545, ZN => n5044);
   U3107 : AOI22_X1 port map( A1 => REGISTERS_16_34_port, A2 => n656, B1 => 
                           REGISTERS_18_34_port, B2 => n619, ZN => n5043);
   U3108 : AND4_X1 port map( A1 => n5046, A2 => n5045, A3 => n5044, A4 => n5043
                           , ZN => n5063);
   U3109 : AOI22_X1 port map( A1 => REGISTERS_29_34_port, A2 => n434, B1 => 
                           REGISTERS_31_34_port, B2 => n397, ZN => n5050);
   U3110 : AOI22_X1 port map( A1 => REGISTERS_25_34_port, A2 => n508, B1 => 
                           REGISTERS_27_34_port, B2 => n471, ZN => n5049);
   U3111 : AOI22_X1 port map( A1 => REGISTERS_28_34_port, A2 => n582, B1 => 
                           REGISTERS_30_34_port, B2 => n545, ZN => n5048);
   U3112 : AOI22_X1 port map( A1 => REGISTERS_24_34_port, A2 => n656, B1 => 
                           REGISTERS_26_34_port, B2 => n619, ZN => n5047);
   U3113 : AND4_X1 port map( A1 => n5050, A2 => n5049, A3 => n5048, A4 => n5047
                           , ZN => n5062);
   U3114 : AOI22_X1 port map( A1 => REGISTERS_5_34_port, A2 => n434, B1 => 
                           REGISTERS_7_34_port, B2 => n397, ZN => n5054);
   U3115 : AOI22_X1 port map( A1 => REGISTERS_1_34_port, A2 => n508, B1 => 
                           REGISTERS_3_34_port, B2 => n471, ZN => n5053);
   U3116 : AOI22_X1 port map( A1 => REGISTERS_4_34_port, A2 => n582, B1 => 
                           REGISTERS_6_34_port, B2 => n545, ZN => n5052);
   U3117 : AOI22_X1 port map( A1 => REGISTERS_0_34_port, A2 => n656, B1 => 
                           REGISTERS_2_34_port, B2 => n619, ZN => n5051);
   U3118 : NAND4_X1 port map( A1 => n5054, A2 => n5053, A3 => n5052, A4 => 
                           n5051, ZN => n5060);
   U3119 : AOI22_X1 port map( A1 => REGISTERS_13_34_port, A2 => n434, B1 => 
                           REGISTERS_15_34_port, B2 => n397, ZN => n5058);
   U3120 : AOI22_X1 port map( A1 => REGISTERS_9_34_port, A2 => n508, B1 => 
                           REGISTERS_11_34_port, B2 => n471, ZN => n5057);
   U3121 : AOI22_X1 port map( A1 => REGISTERS_12_34_port, A2 => n582, B1 => 
                           REGISTERS_14_34_port, B2 => n545, ZN => n5056);
   U3122 : AOI22_X1 port map( A1 => REGISTERS_8_34_port, A2 => n656, B1 => 
                           REGISTERS_10_34_port, B2 => n619, ZN => n5055);
   U3123 : NAND4_X1 port map( A1 => n5058, A2 => n5057, A3 => n5056, A4 => 
                           n5055, ZN => n5059);
   U3124 : AOI22_X1 port map( A1 => n5060, A2 => n23, B1 => n5059, B2 => n22, 
                           ZN => n5061);
   U3125 : OAI221_X1 port map( B1 => n5673, B2 => n5063, C1 => n5671, C2 => 
                           n5062, A => n5061, ZN => N254);
   U3126 : AOI22_X1 port map( A1 => REGISTERS_21_35_port, A2 => n434, B1 => 
                           REGISTERS_23_35_port, B2 => n397, ZN => n5067);
   U3127 : AOI22_X1 port map( A1 => REGISTERS_17_35_port, A2 => n508, B1 => 
                           REGISTERS_19_35_port, B2 => n471, ZN => n5066);
   U3128 : AOI22_X1 port map( A1 => REGISTERS_20_35_port, A2 => n582, B1 => 
                           REGISTERS_22_35_port, B2 => n545, ZN => n5065);
   U3129 : AOI22_X1 port map( A1 => REGISTERS_16_35_port, A2 => n656, B1 => 
                           REGISTERS_18_35_port, B2 => n619, ZN => n5064);
   U3130 : AND4_X1 port map( A1 => n5067, A2 => n5066, A3 => n5065, A4 => n5064
                           , ZN => n5084);
   U3131 : AOI22_X1 port map( A1 => REGISTERS_29_35_port, A2 => n434, B1 => 
                           REGISTERS_31_35_port, B2 => n397, ZN => n5071);
   U3132 : AOI22_X1 port map( A1 => REGISTERS_25_35_port, A2 => n508, B1 => 
                           REGISTERS_27_35_port, B2 => n471, ZN => n5070);
   U3133 : AOI22_X1 port map( A1 => REGISTERS_28_35_port, A2 => n582, B1 => 
                           REGISTERS_30_35_port, B2 => n545, ZN => n5069);
   U3134 : AOI22_X1 port map( A1 => REGISTERS_24_35_port, A2 => n656, B1 => 
                           REGISTERS_26_35_port, B2 => n619, ZN => n5068);
   U3135 : AND4_X1 port map( A1 => n5071, A2 => n5070, A3 => n5069, A4 => n5068
                           , ZN => n5083);
   U3136 : AOI22_X1 port map( A1 => REGISTERS_5_35_port, A2 => n434, B1 => 
                           REGISTERS_7_35_port, B2 => n397, ZN => n5075);
   U3137 : AOI22_X1 port map( A1 => REGISTERS_1_35_port, A2 => n508, B1 => 
                           REGISTERS_3_35_port, B2 => n471, ZN => n5074);
   U3138 : AOI22_X1 port map( A1 => REGISTERS_4_35_port, A2 => n582, B1 => 
                           REGISTERS_6_35_port, B2 => n545, ZN => n5073);
   U3139 : AOI22_X1 port map( A1 => REGISTERS_0_35_port, A2 => n656, B1 => 
                           REGISTERS_2_35_port, B2 => n619, ZN => n5072);
   U3140 : NAND4_X1 port map( A1 => n5075, A2 => n5074, A3 => n5073, A4 => 
                           n5072, ZN => n5081);
   U3141 : AOI22_X1 port map( A1 => REGISTERS_13_35_port, A2 => n434, B1 => 
                           REGISTERS_15_35_port, B2 => n397, ZN => n5079);
   U3142 : AOI22_X1 port map( A1 => REGISTERS_9_35_port, A2 => n508, B1 => 
                           REGISTERS_11_35_port, B2 => n471, ZN => n5078);
   U3143 : AOI22_X1 port map( A1 => REGISTERS_12_35_port, A2 => n582, B1 => 
                           REGISTERS_14_35_port, B2 => n545, ZN => n5077);
   U3144 : AOI22_X1 port map( A1 => REGISTERS_8_35_port, A2 => n656, B1 => 
                           REGISTERS_10_35_port, B2 => n619, ZN => n5076);
   U3145 : NAND4_X1 port map( A1 => n5079, A2 => n5078, A3 => n5077, A4 => 
                           n5076, ZN => n5080);
   U3146 : AOI22_X1 port map( A1 => n5081, A2 => n23, B1 => n5080, B2 => n22, 
                           ZN => n5082);
   U3147 : OAI221_X1 port map( B1 => n5673, B2 => n5084, C1 => n5671, C2 => 
                           n5083, A => n5082, ZN => N253);
   U3148 : AOI22_X1 port map( A1 => REGISTERS_21_36_port, A2 => n435, B1 => 
                           REGISTERS_23_36_port, B2 => n398, ZN => n5088);
   U3149 : AOI22_X1 port map( A1 => REGISTERS_17_36_port, A2 => n509, B1 => 
                           REGISTERS_19_36_port, B2 => n472, ZN => n5087);
   U3150 : AOI22_X1 port map( A1 => REGISTERS_20_36_port, A2 => n583, B1 => 
                           REGISTERS_22_36_port, B2 => n546, ZN => n5086);
   U3151 : AOI22_X1 port map( A1 => REGISTERS_16_36_port, A2 => n657, B1 => 
                           REGISTERS_18_36_port, B2 => n620, ZN => n5085);
   U3152 : AND4_X1 port map( A1 => n5088, A2 => n5087, A3 => n5086, A4 => n5085
                           , ZN => n5105);
   U3153 : AOI22_X1 port map( A1 => REGISTERS_29_36_port, A2 => n435, B1 => 
                           REGISTERS_31_36_port, B2 => n398, ZN => n5092);
   U3154 : AOI22_X1 port map( A1 => REGISTERS_25_36_port, A2 => n509, B1 => 
                           REGISTERS_27_36_port, B2 => n472, ZN => n5091);
   U3155 : AOI22_X1 port map( A1 => REGISTERS_28_36_port, A2 => n583, B1 => 
                           REGISTERS_30_36_port, B2 => n546, ZN => n5090);
   U3156 : AOI22_X1 port map( A1 => REGISTERS_24_36_port, A2 => n657, B1 => 
                           REGISTERS_26_36_port, B2 => n620, ZN => n5089);
   U3157 : AND4_X1 port map( A1 => n5092, A2 => n5091, A3 => n5090, A4 => n5089
                           , ZN => n5104);
   U3158 : AOI22_X1 port map( A1 => REGISTERS_5_36_port, A2 => n435, B1 => 
                           REGISTERS_7_36_port, B2 => n398, ZN => n5096);
   U3159 : AOI22_X1 port map( A1 => REGISTERS_1_36_port, A2 => n509, B1 => 
                           REGISTERS_3_36_port, B2 => n472, ZN => n5095);
   U3160 : AOI22_X1 port map( A1 => REGISTERS_4_36_port, A2 => n583, B1 => 
                           REGISTERS_6_36_port, B2 => n546, ZN => n5094);
   U3161 : AOI22_X1 port map( A1 => REGISTERS_0_36_port, A2 => n657, B1 => 
                           REGISTERS_2_36_port, B2 => n620, ZN => n5093);
   U3162 : NAND4_X1 port map( A1 => n5096, A2 => n5095, A3 => n5094, A4 => 
                           n5093, ZN => n5102);
   U3163 : AOI22_X1 port map( A1 => REGISTERS_13_36_port, A2 => n435, B1 => 
                           REGISTERS_15_36_port, B2 => n398, ZN => n5100);
   U3164 : AOI22_X1 port map( A1 => REGISTERS_9_36_port, A2 => n509, B1 => 
                           REGISTERS_11_36_port, B2 => n472, ZN => n5099);
   U3165 : AOI22_X1 port map( A1 => REGISTERS_12_36_port, A2 => n583, B1 => 
                           REGISTERS_14_36_port, B2 => n546, ZN => n5098);
   U3166 : AOI22_X1 port map( A1 => REGISTERS_8_36_port, A2 => n657, B1 => 
                           REGISTERS_10_36_port, B2 => n620, ZN => n5097);
   U3167 : NAND4_X1 port map( A1 => n5100, A2 => n5099, A3 => n5098, A4 => 
                           n5097, ZN => n5101);
   U3168 : AOI22_X1 port map( A1 => n5102, A2 => n23, B1 => n5101, B2 => n22, 
                           ZN => n5103);
   U3169 : OAI221_X1 port map( B1 => n5673, B2 => n5105, C1 => n5671, C2 => 
                           n5104, A => n5103, ZN => N252);
   U3170 : AOI22_X1 port map( A1 => REGISTERS_21_37_port, A2 => n435, B1 => 
                           REGISTERS_23_37_port, B2 => n398, ZN => n5109);
   U3171 : AOI22_X1 port map( A1 => REGISTERS_17_37_port, A2 => n509, B1 => 
                           REGISTERS_19_37_port, B2 => n472, ZN => n5108);
   U3172 : AOI22_X1 port map( A1 => REGISTERS_20_37_port, A2 => n583, B1 => 
                           REGISTERS_22_37_port, B2 => n546, ZN => n5107);
   U3173 : AOI22_X1 port map( A1 => REGISTERS_16_37_port, A2 => n657, B1 => 
                           REGISTERS_18_37_port, B2 => n620, ZN => n5106);
   U3174 : AND4_X1 port map( A1 => n5109, A2 => n5108, A3 => n5107, A4 => n5106
                           , ZN => n5126);
   U3175 : AOI22_X1 port map( A1 => REGISTERS_29_37_port, A2 => n435, B1 => 
                           REGISTERS_31_37_port, B2 => n398, ZN => n5113);
   U3176 : AOI22_X1 port map( A1 => REGISTERS_25_37_port, A2 => n509, B1 => 
                           REGISTERS_27_37_port, B2 => n472, ZN => n5112);
   U3177 : AOI22_X1 port map( A1 => REGISTERS_28_37_port, A2 => n583, B1 => 
                           REGISTERS_30_37_port, B2 => n546, ZN => n5111);
   U3178 : AOI22_X1 port map( A1 => REGISTERS_24_37_port, A2 => n657, B1 => 
                           REGISTERS_26_37_port, B2 => n620, ZN => n5110);
   U3179 : AND4_X1 port map( A1 => n5113, A2 => n5112, A3 => n5111, A4 => n5110
                           , ZN => n5125);
   U3180 : AOI22_X1 port map( A1 => REGISTERS_5_37_port, A2 => n435, B1 => 
                           REGISTERS_7_37_port, B2 => n398, ZN => n5117);
   U3181 : AOI22_X1 port map( A1 => REGISTERS_1_37_port, A2 => n509, B1 => 
                           REGISTERS_3_37_port, B2 => n472, ZN => n5116);
   U3182 : AOI22_X1 port map( A1 => REGISTERS_4_37_port, A2 => n583, B1 => 
                           REGISTERS_6_37_port, B2 => n546, ZN => n5115);
   U3183 : AOI22_X1 port map( A1 => REGISTERS_0_37_port, A2 => n657, B1 => 
                           REGISTERS_2_37_port, B2 => n620, ZN => n5114);
   U3184 : NAND4_X1 port map( A1 => n5117, A2 => n5116, A3 => n5115, A4 => 
                           n5114, ZN => n5123);
   U3185 : AOI22_X1 port map( A1 => REGISTERS_13_37_port, A2 => n435, B1 => 
                           REGISTERS_15_37_port, B2 => n398, ZN => n5121);
   U3186 : AOI22_X1 port map( A1 => REGISTERS_9_37_port, A2 => n509, B1 => 
                           REGISTERS_11_37_port, B2 => n472, ZN => n5120);
   U3187 : AOI22_X1 port map( A1 => REGISTERS_12_37_port, A2 => n583, B1 => 
                           REGISTERS_14_37_port, B2 => n546, ZN => n5119);
   U3188 : AOI22_X1 port map( A1 => REGISTERS_8_37_port, A2 => n657, B1 => 
                           REGISTERS_10_37_port, B2 => n620, ZN => n5118);
   U3189 : NAND4_X1 port map( A1 => n5121, A2 => n5120, A3 => n5119, A4 => 
                           n5118, ZN => n5122);
   U3190 : AOI22_X1 port map( A1 => n5123, A2 => n23, B1 => n5122, B2 => n22, 
                           ZN => n5124);
   U3191 : OAI221_X1 port map( B1 => n5673, B2 => n5126, C1 => n5671, C2 => 
                           n5125, A => n5124, ZN => N251);
   U3192 : AOI22_X1 port map( A1 => REGISTERS_21_38_port, A2 => n435, B1 => 
                           REGISTERS_23_38_port, B2 => n398, ZN => n5130);
   U3193 : AOI22_X1 port map( A1 => REGISTERS_17_38_port, A2 => n509, B1 => 
                           REGISTERS_19_38_port, B2 => n472, ZN => n5129);
   U3194 : AOI22_X1 port map( A1 => REGISTERS_20_38_port, A2 => n583, B1 => 
                           REGISTERS_22_38_port, B2 => n546, ZN => n5128);
   U3195 : AOI22_X1 port map( A1 => REGISTERS_16_38_port, A2 => n657, B1 => 
                           REGISTERS_18_38_port, B2 => n620, ZN => n5127);
   U3196 : AND4_X1 port map( A1 => n5130, A2 => n5129, A3 => n5128, A4 => n5127
                           , ZN => n5147);
   U3197 : AOI22_X1 port map( A1 => REGISTERS_29_38_port, A2 => n435, B1 => 
                           REGISTERS_31_38_port, B2 => n398, ZN => n5134);
   U3198 : AOI22_X1 port map( A1 => REGISTERS_25_38_port, A2 => n509, B1 => 
                           REGISTERS_27_38_port, B2 => n472, ZN => n5133);
   U3199 : AOI22_X1 port map( A1 => REGISTERS_28_38_port, A2 => n583, B1 => 
                           REGISTERS_30_38_port, B2 => n546, ZN => n5132);
   U3200 : AOI22_X1 port map( A1 => REGISTERS_24_38_port, A2 => n657, B1 => 
                           REGISTERS_26_38_port, B2 => n620, ZN => n5131);
   U3201 : AND4_X1 port map( A1 => n5134, A2 => n5133, A3 => n5132, A4 => n5131
                           , ZN => n5146);
   U3202 : AOI22_X1 port map( A1 => REGISTERS_5_38_port, A2 => n435, B1 => 
                           REGISTERS_7_38_port, B2 => n398, ZN => n5138);
   U3203 : AOI22_X1 port map( A1 => REGISTERS_1_38_port, A2 => n509, B1 => 
                           REGISTERS_3_38_port, B2 => n472, ZN => n5137);
   U3204 : AOI22_X1 port map( A1 => REGISTERS_4_38_port, A2 => n583, B1 => 
                           REGISTERS_6_38_port, B2 => n546, ZN => n5136);
   U3205 : AOI22_X1 port map( A1 => REGISTERS_0_38_port, A2 => n657, B1 => 
                           REGISTERS_2_38_port, B2 => n620, ZN => n5135);
   U3206 : NAND4_X1 port map( A1 => n5138, A2 => n5137, A3 => n5136, A4 => 
                           n5135, ZN => n5144);
   U3207 : AOI22_X1 port map( A1 => REGISTERS_13_38_port, A2 => n435, B1 => 
                           REGISTERS_15_38_port, B2 => n398, ZN => n5142);
   U3208 : AOI22_X1 port map( A1 => REGISTERS_9_38_port, A2 => n509, B1 => 
                           REGISTERS_11_38_port, B2 => n472, ZN => n5141);
   U3209 : AOI22_X1 port map( A1 => REGISTERS_12_38_port, A2 => n583, B1 => 
                           REGISTERS_14_38_port, B2 => n546, ZN => n5140);
   U3210 : AOI22_X1 port map( A1 => REGISTERS_8_38_port, A2 => n657, B1 => 
                           REGISTERS_10_38_port, B2 => n620, ZN => n5139);
   U3211 : NAND4_X1 port map( A1 => n5142, A2 => n5141, A3 => n5140, A4 => 
                           n5139, ZN => n5143);
   U3212 : AOI22_X1 port map( A1 => n5144, A2 => n23, B1 => n5143, B2 => n22, 
                           ZN => n5145);
   U3213 : OAI221_X1 port map( B1 => n5673, B2 => n5147, C1 => n5671, C2 => 
                           n5146, A => n5145, ZN => N250);
   U3214 : AOI22_X1 port map( A1 => REGISTERS_21_39_port, A2 => n436, B1 => 
                           REGISTERS_23_39_port, B2 => n399, ZN => n5151);
   U3215 : AOI22_X1 port map( A1 => REGISTERS_17_39_port, A2 => n510, B1 => 
                           REGISTERS_19_39_port, B2 => n473, ZN => n5150);
   U3216 : AOI22_X1 port map( A1 => REGISTERS_20_39_port, A2 => n584, B1 => 
                           REGISTERS_22_39_port, B2 => n547, ZN => n5149);
   U3217 : AOI22_X1 port map( A1 => REGISTERS_16_39_port, A2 => n658, B1 => 
                           REGISTERS_18_39_port, B2 => n621, ZN => n5148);
   U3218 : AND4_X1 port map( A1 => n5151, A2 => n5150, A3 => n5149, A4 => n5148
                           , ZN => n5168);
   U3219 : AOI22_X1 port map( A1 => REGISTERS_29_39_port, A2 => n436, B1 => 
                           REGISTERS_31_39_port, B2 => n399, ZN => n5155);
   U3220 : AOI22_X1 port map( A1 => REGISTERS_25_39_port, A2 => n510, B1 => 
                           REGISTERS_27_39_port, B2 => n473, ZN => n5154);
   U3221 : AOI22_X1 port map( A1 => REGISTERS_28_39_port, A2 => n584, B1 => 
                           REGISTERS_30_39_port, B2 => n547, ZN => n5153);
   U3222 : AOI22_X1 port map( A1 => REGISTERS_24_39_port, A2 => n658, B1 => 
                           REGISTERS_26_39_port, B2 => n621, ZN => n5152);
   U3223 : AND4_X1 port map( A1 => n5155, A2 => n5154, A3 => n5153, A4 => n5152
                           , ZN => n5167);
   U3224 : AOI22_X1 port map( A1 => REGISTERS_5_39_port, A2 => n436, B1 => 
                           REGISTERS_7_39_port, B2 => n399, ZN => n5159);
   U3225 : AOI22_X1 port map( A1 => REGISTERS_1_39_port, A2 => n510, B1 => 
                           REGISTERS_3_39_port, B2 => n473, ZN => n5158);
   U3226 : AOI22_X1 port map( A1 => REGISTERS_4_39_port, A2 => n584, B1 => 
                           REGISTERS_6_39_port, B2 => n547, ZN => n5157);
   U3227 : AOI22_X1 port map( A1 => REGISTERS_0_39_port, A2 => n658, B1 => 
                           REGISTERS_2_39_port, B2 => n621, ZN => n5156);
   U3228 : NAND4_X1 port map( A1 => n5159, A2 => n5158, A3 => n5157, A4 => 
                           n5156, ZN => n5165);
   U3229 : AOI22_X1 port map( A1 => REGISTERS_13_39_port, A2 => n436, B1 => 
                           REGISTERS_15_39_port, B2 => n399, ZN => n5163);
   U3230 : AOI22_X1 port map( A1 => REGISTERS_9_39_port, A2 => n510, B1 => 
                           REGISTERS_11_39_port, B2 => n473, ZN => n5162);
   U3231 : AOI22_X1 port map( A1 => REGISTERS_12_39_port, A2 => n584, B1 => 
                           REGISTERS_14_39_port, B2 => n547, ZN => n5161);
   U3232 : AOI22_X1 port map( A1 => REGISTERS_8_39_port, A2 => n658, B1 => 
                           REGISTERS_10_39_port, B2 => n621, ZN => n5160);
   U3233 : NAND4_X1 port map( A1 => n5163, A2 => n5162, A3 => n5161, A4 => 
                           n5160, ZN => n5164);
   U3234 : AOI22_X1 port map( A1 => n5165, A2 => n23, B1 => n5164, B2 => n22, 
                           ZN => n5166);
   U3235 : OAI221_X1 port map( B1 => n5673, B2 => n5168, C1 => n5671, C2 => 
                           n5167, A => n5166, ZN => N249);
   U3236 : AOI22_X1 port map( A1 => REGISTERS_21_40_port, A2 => n436, B1 => 
                           REGISTERS_23_40_port, B2 => n399, ZN => n5172);
   U3237 : AOI22_X1 port map( A1 => REGISTERS_17_40_port, A2 => n510, B1 => 
                           REGISTERS_19_40_port, B2 => n473, ZN => n5171);
   U3238 : AOI22_X1 port map( A1 => REGISTERS_20_40_port, A2 => n584, B1 => 
                           REGISTERS_22_40_port, B2 => n547, ZN => n5170);
   U3239 : AOI22_X1 port map( A1 => REGISTERS_16_40_port, A2 => n658, B1 => 
                           REGISTERS_18_40_port, B2 => n621, ZN => n5169);
   U3240 : AND4_X1 port map( A1 => n5172, A2 => n5171, A3 => n5170, A4 => n5169
                           , ZN => n5189);
   U3241 : AOI22_X1 port map( A1 => REGISTERS_29_40_port, A2 => n436, B1 => 
                           REGISTERS_31_40_port, B2 => n399, ZN => n5176);
   U3242 : AOI22_X1 port map( A1 => REGISTERS_25_40_port, A2 => n510, B1 => 
                           REGISTERS_27_40_port, B2 => n473, ZN => n5175);
   U3243 : AOI22_X1 port map( A1 => REGISTERS_28_40_port, A2 => n584, B1 => 
                           REGISTERS_30_40_port, B2 => n547, ZN => n5174);
   U3244 : AOI22_X1 port map( A1 => REGISTERS_24_40_port, A2 => n658, B1 => 
                           REGISTERS_26_40_port, B2 => n621, ZN => n5173);
   U3245 : AND4_X1 port map( A1 => n5176, A2 => n5175, A3 => n5174, A4 => n5173
                           , ZN => n5188);
   U3246 : AOI22_X1 port map( A1 => REGISTERS_5_40_port, A2 => n436, B1 => 
                           REGISTERS_7_40_port, B2 => n399, ZN => n5180);
   U3247 : AOI22_X1 port map( A1 => REGISTERS_1_40_port, A2 => n510, B1 => 
                           REGISTERS_3_40_port, B2 => n473, ZN => n5179);
   U3248 : AOI22_X1 port map( A1 => REGISTERS_4_40_port, A2 => n584, B1 => 
                           REGISTERS_6_40_port, B2 => n547, ZN => n5178);
   U3249 : AOI22_X1 port map( A1 => REGISTERS_0_40_port, A2 => n658, B1 => 
                           REGISTERS_2_40_port, B2 => n621, ZN => n5177);
   U3250 : NAND4_X1 port map( A1 => n5180, A2 => n5179, A3 => n5178, A4 => 
                           n5177, ZN => n5186);
   U3251 : AOI22_X1 port map( A1 => REGISTERS_13_40_port, A2 => n436, B1 => 
                           REGISTERS_15_40_port, B2 => n399, ZN => n5184);
   U3252 : AOI22_X1 port map( A1 => REGISTERS_9_40_port, A2 => n510, B1 => 
                           REGISTERS_11_40_port, B2 => n473, ZN => n5183);
   U3253 : AOI22_X1 port map( A1 => REGISTERS_12_40_port, A2 => n584, B1 => 
                           REGISTERS_14_40_port, B2 => n547, ZN => n5182);
   U3254 : AOI22_X1 port map( A1 => REGISTERS_8_40_port, A2 => n658, B1 => 
                           REGISTERS_10_40_port, B2 => n621, ZN => n5181);
   U3255 : NAND4_X1 port map( A1 => n5184, A2 => n5183, A3 => n5182, A4 => 
                           n5181, ZN => n5185);
   U3256 : AOI22_X1 port map( A1 => n5186, A2 => n23, B1 => n5185, B2 => n22, 
                           ZN => n5187);
   U3257 : OAI221_X1 port map( B1 => n5673, B2 => n5189, C1 => n5671, C2 => 
                           n5188, A => n5187, ZN => N248);
   U3258 : AOI22_X1 port map( A1 => REGISTERS_21_41_port, A2 => n436, B1 => 
                           REGISTERS_23_41_port, B2 => n399, ZN => n5193);
   U3259 : AOI22_X1 port map( A1 => REGISTERS_17_41_port, A2 => n510, B1 => 
                           REGISTERS_19_41_port, B2 => n473, ZN => n5192);
   U3260 : AOI22_X1 port map( A1 => REGISTERS_20_41_port, A2 => n584, B1 => 
                           REGISTERS_22_41_port, B2 => n547, ZN => n5191);
   U3261 : AOI22_X1 port map( A1 => REGISTERS_16_41_port, A2 => n658, B1 => 
                           REGISTERS_18_41_port, B2 => n621, ZN => n5190);
   U3262 : AND4_X1 port map( A1 => n5193, A2 => n5192, A3 => n5191, A4 => n5190
                           , ZN => n5210);
   U3263 : AOI22_X1 port map( A1 => REGISTERS_29_41_port, A2 => n436, B1 => 
                           REGISTERS_31_41_port, B2 => n399, ZN => n5197);
   U3264 : AOI22_X1 port map( A1 => REGISTERS_25_41_port, A2 => n510, B1 => 
                           REGISTERS_27_41_port, B2 => n473, ZN => n5196);
   U3265 : AOI22_X1 port map( A1 => REGISTERS_28_41_port, A2 => n584, B1 => 
                           REGISTERS_30_41_port, B2 => n547, ZN => n5195);
   U3266 : AOI22_X1 port map( A1 => REGISTERS_24_41_port, A2 => n658, B1 => 
                           REGISTERS_26_41_port, B2 => n621, ZN => n5194);
   U3267 : AND4_X1 port map( A1 => n5197, A2 => n5196, A3 => n5195, A4 => n5194
                           , ZN => n5209);
   U3268 : AOI22_X1 port map( A1 => REGISTERS_5_41_port, A2 => n436, B1 => 
                           REGISTERS_7_41_port, B2 => n399, ZN => n5201);
   U3269 : AOI22_X1 port map( A1 => REGISTERS_1_41_port, A2 => n510, B1 => 
                           REGISTERS_3_41_port, B2 => n473, ZN => n5200);
   U3270 : AOI22_X1 port map( A1 => REGISTERS_4_41_port, A2 => n584, B1 => 
                           REGISTERS_6_41_port, B2 => n547, ZN => n5199);
   U3271 : AOI22_X1 port map( A1 => REGISTERS_0_41_port, A2 => n658, B1 => 
                           REGISTERS_2_41_port, B2 => n621, ZN => n5198);
   U3272 : NAND4_X1 port map( A1 => n5201, A2 => n5200, A3 => n5199, A4 => 
                           n5198, ZN => n5207);
   U3273 : AOI22_X1 port map( A1 => REGISTERS_13_41_port, A2 => n436, B1 => 
                           REGISTERS_15_41_port, B2 => n399, ZN => n5205);
   U3274 : AOI22_X1 port map( A1 => REGISTERS_9_41_port, A2 => n510, B1 => 
                           REGISTERS_11_41_port, B2 => n473, ZN => n5204);
   U3275 : AOI22_X1 port map( A1 => REGISTERS_12_41_port, A2 => n584, B1 => 
                           REGISTERS_14_41_port, B2 => n547, ZN => n5203);
   U3276 : AOI22_X1 port map( A1 => REGISTERS_8_41_port, A2 => n658, B1 => 
                           REGISTERS_10_41_port, B2 => n621, ZN => n5202);
   U3277 : NAND4_X1 port map( A1 => n5205, A2 => n5204, A3 => n5203, A4 => 
                           n5202, ZN => n5206);
   U3278 : AOI22_X1 port map( A1 => n5207, A2 => n23, B1 => n5206, B2 => n22, 
                           ZN => n5208);
   U3279 : OAI221_X1 port map( B1 => n5673, B2 => n5210, C1 => n5671, C2 => 
                           n5209, A => n5208, ZN => N247);
   U3280 : AOI22_X1 port map( A1 => REGISTERS_21_42_port, A2 => n437, B1 => 
                           REGISTERS_23_42_port, B2 => n400, ZN => n5214);
   U3281 : AOI22_X1 port map( A1 => REGISTERS_17_42_port, A2 => n511, B1 => 
                           REGISTERS_19_42_port, B2 => n474, ZN => n5213);
   U3282 : AOI22_X1 port map( A1 => REGISTERS_20_42_port, A2 => n585, B1 => 
                           REGISTERS_22_42_port, B2 => n548, ZN => n5212);
   U3283 : AOI22_X1 port map( A1 => REGISTERS_16_42_port, A2 => n659, B1 => 
                           REGISTERS_18_42_port, B2 => n622, ZN => n5211);
   U3284 : AND4_X1 port map( A1 => n5214, A2 => n5213, A3 => n5212, A4 => n5211
                           , ZN => n5231);
   U3285 : AOI22_X1 port map( A1 => REGISTERS_29_42_port, A2 => n437, B1 => 
                           REGISTERS_31_42_port, B2 => n400, ZN => n5218);
   U3286 : AOI22_X1 port map( A1 => REGISTERS_25_42_port, A2 => n511, B1 => 
                           REGISTERS_27_42_port, B2 => n474, ZN => n5217);
   U3287 : AOI22_X1 port map( A1 => REGISTERS_28_42_port, A2 => n585, B1 => 
                           REGISTERS_30_42_port, B2 => n548, ZN => n5216);
   U3288 : AOI22_X1 port map( A1 => REGISTERS_24_42_port, A2 => n659, B1 => 
                           REGISTERS_26_42_port, B2 => n622, ZN => n5215);
   U3289 : AND4_X1 port map( A1 => n5218, A2 => n5217, A3 => n5216, A4 => n5215
                           , ZN => n5230);
   U3290 : AOI22_X1 port map( A1 => REGISTERS_5_42_port, A2 => n437, B1 => 
                           REGISTERS_7_42_port, B2 => n400, ZN => n5222);
   U3291 : AOI22_X1 port map( A1 => REGISTERS_1_42_port, A2 => n511, B1 => 
                           REGISTERS_3_42_port, B2 => n474, ZN => n5221);
   U3292 : AOI22_X1 port map( A1 => REGISTERS_4_42_port, A2 => n585, B1 => 
                           REGISTERS_6_42_port, B2 => n548, ZN => n5220);
   U3293 : AOI22_X1 port map( A1 => REGISTERS_0_42_port, A2 => n659, B1 => 
                           REGISTERS_2_42_port, B2 => n622, ZN => n5219);
   U3294 : NAND4_X1 port map( A1 => n5222, A2 => n5221, A3 => n5220, A4 => 
                           n5219, ZN => n5228);
   U3295 : AOI22_X1 port map( A1 => REGISTERS_13_42_port, A2 => n437, B1 => 
                           REGISTERS_15_42_port, B2 => n400, ZN => n5226);
   U3296 : AOI22_X1 port map( A1 => REGISTERS_9_42_port, A2 => n511, B1 => 
                           REGISTERS_11_42_port, B2 => n474, ZN => n5225);
   U3297 : AOI22_X1 port map( A1 => REGISTERS_12_42_port, A2 => n585, B1 => 
                           REGISTERS_14_42_port, B2 => n548, ZN => n5224);
   U3298 : AOI22_X1 port map( A1 => REGISTERS_8_42_port, A2 => n659, B1 => 
                           REGISTERS_10_42_port, B2 => n622, ZN => n5223);
   U3299 : NAND4_X1 port map( A1 => n5226, A2 => n5225, A3 => n5224, A4 => 
                           n5223, ZN => n5227);
   U3300 : AOI22_X1 port map( A1 => n5228, A2 => n23, B1 => n5227, B2 => n22, 
                           ZN => n5229);
   U3301 : OAI221_X1 port map( B1 => n5673, B2 => n5231, C1 => n5671, C2 => 
                           n5230, A => n5229, ZN => N246);
   U3302 : AOI22_X1 port map( A1 => REGISTERS_21_43_port, A2 => n437, B1 => 
                           REGISTERS_23_43_port, B2 => n400, ZN => n5235);
   U3303 : AOI22_X1 port map( A1 => REGISTERS_17_43_port, A2 => n511, B1 => 
                           REGISTERS_19_43_port, B2 => n474, ZN => n5234);
   U3304 : AOI22_X1 port map( A1 => REGISTERS_20_43_port, A2 => n585, B1 => 
                           REGISTERS_22_43_port, B2 => n548, ZN => n5233);
   U3305 : AOI22_X1 port map( A1 => REGISTERS_16_43_port, A2 => n659, B1 => 
                           REGISTERS_18_43_port, B2 => n622, ZN => n5232);
   U3306 : AND4_X1 port map( A1 => n5235, A2 => n5234, A3 => n5233, A4 => n5232
                           , ZN => n5252);
   U3307 : AOI22_X1 port map( A1 => REGISTERS_29_43_port, A2 => n437, B1 => 
                           REGISTERS_31_43_port, B2 => n400, ZN => n5239);
   U3308 : AOI22_X1 port map( A1 => REGISTERS_25_43_port, A2 => n511, B1 => 
                           REGISTERS_27_43_port, B2 => n474, ZN => n5238);
   U3309 : AOI22_X1 port map( A1 => REGISTERS_28_43_port, A2 => n585, B1 => 
                           REGISTERS_30_43_port, B2 => n548, ZN => n5237);
   U3310 : AOI22_X1 port map( A1 => REGISTERS_24_43_port, A2 => n659, B1 => 
                           REGISTERS_26_43_port, B2 => n622, ZN => n5236);
   U3311 : AND4_X1 port map( A1 => n5239, A2 => n5238, A3 => n5237, A4 => n5236
                           , ZN => n5251);
   U3312 : AOI22_X1 port map( A1 => REGISTERS_5_43_port, A2 => n437, B1 => 
                           REGISTERS_7_43_port, B2 => n400, ZN => n5243);
   U3313 : AOI22_X1 port map( A1 => REGISTERS_1_43_port, A2 => n511, B1 => 
                           REGISTERS_3_43_port, B2 => n474, ZN => n5242);
   U3314 : AOI22_X1 port map( A1 => REGISTERS_4_43_port, A2 => n585, B1 => 
                           REGISTERS_6_43_port, B2 => n548, ZN => n5241);
   U3315 : AOI22_X1 port map( A1 => REGISTERS_0_43_port, A2 => n659, B1 => 
                           REGISTERS_2_43_port, B2 => n622, ZN => n5240);
   U3316 : NAND4_X1 port map( A1 => n5243, A2 => n5242, A3 => n5241, A4 => 
                           n5240, ZN => n5249);
   U3317 : AOI22_X1 port map( A1 => REGISTERS_13_43_port, A2 => n437, B1 => 
                           REGISTERS_15_43_port, B2 => n400, ZN => n5247);
   U3318 : AOI22_X1 port map( A1 => REGISTERS_9_43_port, A2 => n511, B1 => 
                           REGISTERS_11_43_port, B2 => n474, ZN => n5246);
   U3319 : AOI22_X1 port map( A1 => REGISTERS_12_43_port, A2 => n585, B1 => 
                           REGISTERS_14_43_port, B2 => n548, ZN => n5245);
   U3320 : AOI22_X1 port map( A1 => REGISTERS_8_43_port, A2 => n659, B1 => 
                           REGISTERS_10_43_port, B2 => n622, ZN => n5244);
   U3321 : NAND4_X1 port map( A1 => n5247, A2 => n5246, A3 => n5245, A4 => 
                           n5244, ZN => n5248);
   U3322 : AOI22_X1 port map( A1 => n5249, A2 => n23, B1 => n5248, B2 => n22, 
                           ZN => n5250);
   U3323 : OAI221_X1 port map( B1 => n5673, B2 => n5252, C1 => n5671, C2 => 
                           n5251, A => n5250, ZN => N245);
   U3324 : AOI22_X1 port map( A1 => REGISTERS_21_44_port, A2 => n437, B1 => 
                           REGISTERS_23_44_port, B2 => n400, ZN => n5256);
   U3325 : AOI22_X1 port map( A1 => REGISTERS_17_44_port, A2 => n511, B1 => 
                           REGISTERS_19_44_port, B2 => n474, ZN => n5255);
   U3326 : AOI22_X1 port map( A1 => REGISTERS_20_44_port, A2 => n585, B1 => 
                           REGISTERS_22_44_port, B2 => n548, ZN => n5254);
   U3327 : AOI22_X1 port map( A1 => REGISTERS_16_44_port, A2 => n659, B1 => 
                           REGISTERS_18_44_port, B2 => n622, ZN => n5253);
   U3328 : AND4_X1 port map( A1 => n5256, A2 => n5255, A3 => n5254, A4 => n5253
                           , ZN => n5273);
   U3329 : AOI22_X1 port map( A1 => REGISTERS_29_44_port, A2 => n437, B1 => 
                           REGISTERS_31_44_port, B2 => n400, ZN => n5260);
   U3330 : AOI22_X1 port map( A1 => REGISTERS_25_44_port, A2 => n511, B1 => 
                           REGISTERS_27_44_port, B2 => n474, ZN => n5259);
   U3331 : AOI22_X1 port map( A1 => REGISTERS_28_44_port, A2 => n585, B1 => 
                           REGISTERS_30_44_port, B2 => n548, ZN => n5258);
   U3332 : AOI22_X1 port map( A1 => REGISTERS_24_44_port, A2 => n659, B1 => 
                           REGISTERS_26_44_port, B2 => n622, ZN => n5257);
   U3333 : AND4_X1 port map( A1 => n5260, A2 => n5259, A3 => n5258, A4 => n5257
                           , ZN => n5272);
   U3334 : AOI22_X1 port map( A1 => REGISTERS_5_44_port, A2 => n437, B1 => 
                           REGISTERS_7_44_port, B2 => n400, ZN => n5264);
   U3335 : AOI22_X1 port map( A1 => REGISTERS_1_44_port, A2 => n511, B1 => 
                           REGISTERS_3_44_port, B2 => n474, ZN => n5263);
   U3336 : AOI22_X1 port map( A1 => REGISTERS_4_44_port, A2 => n585, B1 => 
                           REGISTERS_6_44_port, B2 => n548, ZN => n5262);
   U3337 : AOI22_X1 port map( A1 => REGISTERS_0_44_port, A2 => n659, B1 => 
                           REGISTERS_2_44_port, B2 => n622, ZN => n5261);
   U3338 : NAND4_X1 port map( A1 => n5264, A2 => n5263, A3 => n5262, A4 => 
                           n5261, ZN => n5270);
   U3339 : AOI22_X1 port map( A1 => REGISTERS_13_44_port, A2 => n437, B1 => 
                           REGISTERS_15_44_port, B2 => n400, ZN => n5268);
   U3340 : AOI22_X1 port map( A1 => REGISTERS_9_44_port, A2 => n511, B1 => 
                           REGISTERS_11_44_port, B2 => n474, ZN => n5267);
   U3341 : AOI22_X1 port map( A1 => REGISTERS_12_44_port, A2 => n585, B1 => 
                           REGISTERS_14_44_port, B2 => n548, ZN => n5266);
   U3342 : AOI22_X1 port map( A1 => REGISTERS_8_44_port, A2 => n659, B1 => 
                           REGISTERS_10_44_port, B2 => n622, ZN => n5265);
   U3343 : NAND4_X1 port map( A1 => n5268, A2 => n5267, A3 => n5266, A4 => 
                           n5265, ZN => n5269);
   U3344 : AOI22_X1 port map( A1 => n5270, A2 => n23, B1 => n5269, B2 => n22, 
                           ZN => n5271);
   U3345 : OAI221_X1 port map( B1 => n5673, B2 => n5273, C1 => n5671, C2 => 
                           n5272, A => n5271, ZN => N244);
   U3346 : AOI22_X1 port map( A1 => REGISTERS_21_45_port, A2 => n438, B1 => 
                           REGISTERS_23_45_port, B2 => n401, ZN => n5277);
   U3347 : AOI22_X1 port map( A1 => REGISTERS_17_45_port, A2 => n512, B1 => 
                           REGISTERS_19_45_port, B2 => n475, ZN => n5276);
   U3348 : AOI22_X1 port map( A1 => REGISTERS_20_45_port, A2 => n586, B1 => 
                           REGISTERS_22_45_port, B2 => n549, ZN => n5275);
   U3349 : AOI22_X1 port map( A1 => REGISTERS_16_45_port, A2 => n660, B1 => 
                           REGISTERS_18_45_port, B2 => n623, ZN => n5274);
   U3350 : AND4_X1 port map( A1 => n5277, A2 => n5276, A3 => n5275, A4 => n5274
                           , ZN => n5294);
   U3351 : AOI22_X1 port map( A1 => REGISTERS_29_45_port, A2 => n438, B1 => 
                           REGISTERS_31_45_port, B2 => n401, ZN => n5281);
   U3352 : AOI22_X1 port map( A1 => REGISTERS_25_45_port, A2 => n512, B1 => 
                           REGISTERS_27_45_port, B2 => n475, ZN => n5280);
   U3353 : AOI22_X1 port map( A1 => REGISTERS_28_45_port, A2 => n586, B1 => 
                           REGISTERS_30_45_port, B2 => n549, ZN => n5279);
   U3354 : AOI22_X1 port map( A1 => REGISTERS_24_45_port, A2 => n660, B1 => 
                           REGISTERS_26_45_port, B2 => n623, ZN => n5278);
   U3355 : AND4_X1 port map( A1 => n5281, A2 => n5280, A3 => n5279, A4 => n5278
                           , ZN => n5293);
   U3356 : AOI22_X1 port map( A1 => REGISTERS_5_45_port, A2 => n438, B1 => 
                           REGISTERS_7_45_port, B2 => n401, ZN => n5285);
   U3357 : AOI22_X1 port map( A1 => REGISTERS_1_45_port, A2 => n512, B1 => 
                           REGISTERS_3_45_port, B2 => n475, ZN => n5284);
   U3358 : AOI22_X1 port map( A1 => REGISTERS_4_45_port, A2 => n586, B1 => 
                           REGISTERS_6_45_port, B2 => n549, ZN => n5283);
   U3359 : AOI22_X1 port map( A1 => REGISTERS_0_45_port, A2 => n660, B1 => 
                           REGISTERS_2_45_port, B2 => n623, ZN => n5282);
   U3360 : NAND4_X1 port map( A1 => n5285, A2 => n5284, A3 => n5283, A4 => 
                           n5282, ZN => n5291);
   U3361 : AOI22_X1 port map( A1 => REGISTERS_13_45_port, A2 => n438, B1 => 
                           REGISTERS_15_45_port, B2 => n401, ZN => n5289);
   U3362 : AOI22_X1 port map( A1 => REGISTERS_9_45_port, A2 => n512, B1 => 
                           REGISTERS_11_45_port, B2 => n475, ZN => n5288);
   U3363 : AOI22_X1 port map( A1 => REGISTERS_12_45_port, A2 => n586, B1 => 
                           REGISTERS_14_45_port, B2 => n549, ZN => n5287);
   U3364 : AOI22_X1 port map( A1 => REGISTERS_8_45_port, A2 => n660, B1 => 
                           REGISTERS_10_45_port, B2 => n623, ZN => n5286);
   U3365 : NAND4_X1 port map( A1 => n5289, A2 => n5288, A3 => n5287, A4 => 
                           n5286, ZN => n5290);
   U3366 : AOI22_X1 port map( A1 => n5291, A2 => n23, B1 => n5290, B2 => n22, 
                           ZN => n5292);
   U3367 : OAI221_X1 port map( B1 => n5673, B2 => n5294, C1 => n5671, C2 => 
                           n5293, A => n5292, ZN => N243);
   U3368 : AOI22_X1 port map( A1 => REGISTERS_21_46_port, A2 => n438, B1 => 
                           REGISTERS_23_46_port, B2 => n401, ZN => n5298);
   U3369 : AOI22_X1 port map( A1 => REGISTERS_17_46_port, A2 => n512, B1 => 
                           REGISTERS_19_46_port, B2 => n475, ZN => n5297);
   U3370 : AOI22_X1 port map( A1 => REGISTERS_20_46_port, A2 => n586, B1 => 
                           REGISTERS_22_46_port, B2 => n549, ZN => n5296);
   U3371 : AOI22_X1 port map( A1 => REGISTERS_16_46_port, A2 => n660, B1 => 
                           REGISTERS_18_46_port, B2 => n623, ZN => n5295);
   U3372 : AND4_X1 port map( A1 => n5298, A2 => n5297, A3 => n5296, A4 => n5295
                           , ZN => n5315);
   U3373 : AOI22_X1 port map( A1 => REGISTERS_29_46_port, A2 => n438, B1 => 
                           REGISTERS_31_46_port, B2 => n401, ZN => n5302);
   U3374 : AOI22_X1 port map( A1 => REGISTERS_25_46_port, A2 => n512, B1 => 
                           REGISTERS_27_46_port, B2 => n475, ZN => n5301);
   U3375 : AOI22_X1 port map( A1 => REGISTERS_28_46_port, A2 => n586, B1 => 
                           REGISTERS_30_46_port, B2 => n549, ZN => n5300);
   U3376 : AOI22_X1 port map( A1 => REGISTERS_24_46_port, A2 => n660, B1 => 
                           REGISTERS_26_46_port, B2 => n623, ZN => n5299);
   U3377 : AND4_X1 port map( A1 => n5302, A2 => n5301, A3 => n5300, A4 => n5299
                           , ZN => n5314);
   U3378 : AOI22_X1 port map( A1 => REGISTERS_5_46_port, A2 => n438, B1 => 
                           REGISTERS_7_46_port, B2 => n401, ZN => n5306);
   U3379 : AOI22_X1 port map( A1 => REGISTERS_1_46_port, A2 => n512, B1 => 
                           REGISTERS_3_46_port, B2 => n475, ZN => n5305);
   U3380 : AOI22_X1 port map( A1 => REGISTERS_4_46_port, A2 => n586, B1 => 
                           REGISTERS_6_46_port, B2 => n549, ZN => n5304);
   U3381 : AOI22_X1 port map( A1 => REGISTERS_0_46_port, A2 => n660, B1 => 
                           REGISTERS_2_46_port, B2 => n623, ZN => n5303);
   U3382 : NAND4_X1 port map( A1 => n5306, A2 => n5305, A3 => n5304, A4 => 
                           n5303, ZN => n5312);
   U3383 : AOI22_X1 port map( A1 => REGISTERS_13_46_port, A2 => n438, B1 => 
                           REGISTERS_15_46_port, B2 => n401, ZN => n5310);
   U3384 : AOI22_X1 port map( A1 => REGISTERS_9_46_port, A2 => n512, B1 => 
                           REGISTERS_11_46_port, B2 => n475, ZN => n5309);
   U3385 : AOI22_X1 port map( A1 => REGISTERS_12_46_port, A2 => n586, B1 => 
                           REGISTERS_14_46_port, B2 => n549, ZN => n5308);
   U3386 : AOI22_X1 port map( A1 => REGISTERS_8_46_port, A2 => n660, B1 => 
                           REGISTERS_10_46_port, B2 => n623, ZN => n5307);
   U3387 : NAND4_X1 port map( A1 => n5310, A2 => n5309, A3 => n5308, A4 => 
                           n5307, ZN => n5311);
   U3388 : AOI22_X1 port map( A1 => n5312, A2 => n23, B1 => n5311, B2 => n22, 
                           ZN => n5313);
   U3389 : OAI221_X1 port map( B1 => n5673, B2 => n5315, C1 => n5671, C2 => 
                           n5314, A => n5313, ZN => N242);
   U3390 : AOI22_X1 port map( A1 => REGISTERS_21_47_port, A2 => n438, B1 => 
                           REGISTERS_23_47_port, B2 => n401, ZN => n5319);
   U3391 : AOI22_X1 port map( A1 => REGISTERS_17_47_port, A2 => n512, B1 => 
                           REGISTERS_19_47_port, B2 => n475, ZN => n5318);
   U3392 : AOI22_X1 port map( A1 => REGISTERS_20_47_port, A2 => n586, B1 => 
                           REGISTERS_22_47_port, B2 => n549, ZN => n5317);
   U3393 : AOI22_X1 port map( A1 => REGISTERS_16_47_port, A2 => n660, B1 => 
                           REGISTERS_18_47_port, B2 => n623, ZN => n5316);
   U3394 : AND4_X1 port map( A1 => n5319, A2 => n5318, A3 => n5317, A4 => n5316
                           , ZN => n5336);
   U3395 : AOI22_X1 port map( A1 => REGISTERS_29_47_port, A2 => n438, B1 => 
                           REGISTERS_31_47_port, B2 => n401, ZN => n5323);
   U3396 : AOI22_X1 port map( A1 => REGISTERS_25_47_port, A2 => n512, B1 => 
                           REGISTERS_27_47_port, B2 => n475, ZN => n5322);
   U3397 : AOI22_X1 port map( A1 => REGISTERS_28_47_port, A2 => n586, B1 => 
                           REGISTERS_30_47_port, B2 => n549, ZN => n5321);
   U3398 : AOI22_X1 port map( A1 => REGISTERS_24_47_port, A2 => n660, B1 => 
                           REGISTERS_26_47_port, B2 => n623, ZN => n5320);
   U3399 : AND4_X1 port map( A1 => n5323, A2 => n5322, A3 => n5321, A4 => n5320
                           , ZN => n5335);
   U3400 : AOI22_X1 port map( A1 => REGISTERS_5_47_port, A2 => n438, B1 => 
                           REGISTERS_7_47_port, B2 => n401, ZN => n5327);
   U3401 : AOI22_X1 port map( A1 => REGISTERS_1_47_port, A2 => n512, B1 => 
                           REGISTERS_3_47_port, B2 => n475, ZN => n5326);
   U3402 : AOI22_X1 port map( A1 => REGISTERS_4_47_port, A2 => n586, B1 => 
                           REGISTERS_6_47_port, B2 => n549, ZN => n5325);
   U3403 : AOI22_X1 port map( A1 => REGISTERS_0_47_port, A2 => n660, B1 => 
                           REGISTERS_2_47_port, B2 => n623, ZN => n5324);
   U3404 : NAND4_X1 port map( A1 => n5327, A2 => n5326, A3 => n5325, A4 => 
                           n5324, ZN => n5333);
   U3405 : AOI22_X1 port map( A1 => REGISTERS_13_47_port, A2 => n438, B1 => 
                           REGISTERS_15_47_port, B2 => n401, ZN => n5331);
   U3406 : AOI22_X1 port map( A1 => REGISTERS_9_47_port, A2 => n512, B1 => 
                           REGISTERS_11_47_port, B2 => n475, ZN => n5330);
   U3407 : AOI22_X1 port map( A1 => REGISTERS_12_47_port, A2 => n586, B1 => 
                           REGISTERS_14_47_port, B2 => n549, ZN => n5329);
   U3408 : AOI22_X1 port map( A1 => REGISTERS_8_47_port, A2 => n660, B1 => 
                           REGISTERS_10_47_port, B2 => n623, ZN => n5328);
   U3409 : NAND4_X1 port map( A1 => n5331, A2 => n5330, A3 => n5329, A4 => 
                           n5328, ZN => n5332);
   U3410 : AOI22_X1 port map( A1 => n5333, A2 => n23, B1 => n5332, B2 => n22, 
                           ZN => n5334);
   U3411 : OAI221_X1 port map( B1 => n5673, B2 => n5336, C1 => n5671, C2 => 
                           n5335, A => n5334, ZN => N241);
   U3412 : AOI22_X1 port map( A1 => REGISTERS_21_48_port, A2 => n439, B1 => 
                           REGISTERS_23_48_port, B2 => n402, ZN => n5340);
   U3413 : AOI22_X1 port map( A1 => REGISTERS_17_48_port, A2 => n513, B1 => 
                           REGISTERS_19_48_port, B2 => n476, ZN => n5339);
   U3414 : AOI22_X1 port map( A1 => REGISTERS_20_48_port, A2 => n587, B1 => 
                           REGISTERS_22_48_port, B2 => n550, ZN => n5338);
   U3415 : AOI22_X1 port map( A1 => REGISTERS_16_48_port, A2 => n661, B1 => 
                           REGISTERS_18_48_port, B2 => n624, ZN => n5337);
   U3416 : AND4_X1 port map( A1 => n5340, A2 => n5339, A3 => n5338, A4 => n5337
                           , ZN => n5357);
   U3417 : AOI22_X1 port map( A1 => REGISTERS_29_48_port, A2 => n439, B1 => 
                           REGISTERS_31_48_port, B2 => n402, ZN => n5344);
   U3418 : AOI22_X1 port map( A1 => REGISTERS_25_48_port, A2 => n513, B1 => 
                           REGISTERS_27_48_port, B2 => n476, ZN => n5343);
   U3419 : AOI22_X1 port map( A1 => REGISTERS_28_48_port, A2 => n587, B1 => 
                           REGISTERS_30_48_port, B2 => n550, ZN => n5342);
   U3420 : AOI22_X1 port map( A1 => REGISTERS_24_48_port, A2 => n661, B1 => 
                           REGISTERS_26_48_port, B2 => n624, ZN => n5341);
   U3421 : AND4_X1 port map( A1 => n5344, A2 => n5343, A3 => n5342, A4 => n5341
                           , ZN => n5356);
   U3422 : AOI22_X1 port map( A1 => REGISTERS_5_48_port, A2 => n439, B1 => 
                           REGISTERS_7_48_port, B2 => n402, ZN => n5348);
   U3423 : AOI22_X1 port map( A1 => REGISTERS_1_48_port, A2 => n513, B1 => 
                           REGISTERS_3_48_port, B2 => n476, ZN => n5347);
   U3424 : AOI22_X1 port map( A1 => REGISTERS_4_48_port, A2 => n587, B1 => 
                           REGISTERS_6_48_port, B2 => n550, ZN => n5346);
   U3425 : AOI22_X1 port map( A1 => REGISTERS_0_48_port, A2 => n661, B1 => 
                           REGISTERS_2_48_port, B2 => n624, ZN => n5345);
   U3426 : NAND4_X1 port map( A1 => n5348, A2 => n5347, A3 => n5346, A4 => 
                           n5345, ZN => n5354);
   U3427 : AOI22_X1 port map( A1 => REGISTERS_13_48_port, A2 => n439, B1 => 
                           REGISTERS_15_48_port, B2 => n402, ZN => n5352);
   U3428 : AOI22_X1 port map( A1 => REGISTERS_9_48_port, A2 => n513, B1 => 
                           REGISTERS_11_48_port, B2 => n476, ZN => n5351);
   U3429 : AOI22_X1 port map( A1 => REGISTERS_12_48_port, A2 => n587, B1 => 
                           REGISTERS_14_48_port, B2 => n550, ZN => n5350);
   U3430 : AOI22_X1 port map( A1 => REGISTERS_8_48_port, A2 => n661, B1 => 
                           REGISTERS_10_48_port, B2 => n624, ZN => n5349);
   U3431 : NAND4_X1 port map( A1 => n5352, A2 => n5351, A3 => n5350, A4 => 
                           n5349, ZN => n5353);
   U3432 : AOI22_X1 port map( A1 => n5354, A2 => n23, B1 => n5353, B2 => n22, 
                           ZN => n5355);
   U3433 : OAI221_X1 port map( B1 => n5673, B2 => n5357, C1 => n5671, C2 => 
                           n5356, A => n5355, ZN => N240);
   U3434 : AOI22_X1 port map( A1 => REGISTERS_21_49_port, A2 => n439, B1 => 
                           REGISTERS_23_49_port, B2 => n402, ZN => n5361);
   U3435 : AOI22_X1 port map( A1 => REGISTERS_17_49_port, A2 => n513, B1 => 
                           REGISTERS_19_49_port, B2 => n476, ZN => n5360);
   U3436 : AOI22_X1 port map( A1 => REGISTERS_20_49_port, A2 => n587, B1 => 
                           REGISTERS_22_49_port, B2 => n550, ZN => n5359);
   U3437 : AOI22_X1 port map( A1 => REGISTERS_16_49_port, A2 => n661, B1 => 
                           REGISTERS_18_49_port, B2 => n624, ZN => n5358);
   U3438 : AND4_X1 port map( A1 => n5361, A2 => n5360, A3 => n5359, A4 => n5358
                           , ZN => n5378);
   U3439 : AOI22_X1 port map( A1 => REGISTERS_29_49_port, A2 => n439, B1 => 
                           REGISTERS_31_49_port, B2 => n402, ZN => n5365);
   U3440 : AOI22_X1 port map( A1 => REGISTERS_25_49_port, A2 => n513, B1 => 
                           REGISTERS_27_49_port, B2 => n476, ZN => n5364);
   U3441 : AOI22_X1 port map( A1 => REGISTERS_28_49_port, A2 => n587, B1 => 
                           REGISTERS_30_49_port, B2 => n550, ZN => n5363);
   U3442 : AOI22_X1 port map( A1 => REGISTERS_24_49_port, A2 => n661, B1 => 
                           REGISTERS_26_49_port, B2 => n624, ZN => n5362);
   U3443 : AND4_X1 port map( A1 => n5365, A2 => n5364, A3 => n5363, A4 => n5362
                           , ZN => n5377);
   U3444 : AOI22_X1 port map( A1 => REGISTERS_5_49_port, A2 => n439, B1 => 
                           REGISTERS_7_49_port, B2 => n402, ZN => n5369);
   U3445 : AOI22_X1 port map( A1 => REGISTERS_1_49_port, A2 => n513, B1 => 
                           REGISTERS_3_49_port, B2 => n476, ZN => n5368);
   U3446 : AOI22_X1 port map( A1 => REGISTERS_4_49_port, A2 => n587, B1 => 
                           REGISTERS_6_49_port, B2 => n550, ZN => n5367);
   U3447 : AOI22_X1 port map( A1 => REGISTERS_0_49_port, A2 => n661, B1 => 
                           REGISTERS_2_49_port, B2 => n624, ZN => n5366);
   U3448 : NAND4_X1 port map( A1 => n5369, A2 => n5368, A3 => n5367, A4 => 
                           n5366, ZN => n5375);
   U3449 : AOI22_X1 port map( A1 => REGISTERS_13_49_port, A2 => n439, B1 => 
                           REGISTERS_15_49_port, B2 => n402, ZN => n5373);
   U3450 : AOI22_X1 port map( A1 => REGISTERS_9_49_port, A2 => n513, B1 => 
                           REGISTERS_11_49_port, B2 => n476, ZN => n5372);
   U3451 : AOI22_X1 port map( A1 => REGISTERS_12_49_port, A2 => n587, B1 => 
                           REGISTERS_14_49_port, B2 => n550, ZN => n5371);
   U3452 : AOI22_X1 port map( A1 => REGISTERS_8_49_port, A2 => n661, B1 => 
                           REGISTERS_10_49_port, B2 => n624, ZN => n5370);
   U3453 : NAND4_X1 port map( A1 => n5373, A2 => n5372, A3 => n5371, A4 => 
                           n5370, ZN => n5374);
   U3454 : AOI22_X1 port map( A1 => n5375, A2 => n23, B1 => n5374, B2 => n22, 
                           ZN => n5376);
   U3455 : OAI221_X1 port map( B1 => n5673, B2 => n5378, C1 => n5671, C2 => 
                           n5377, A => n5376, ZN => N239);
   U3456 : AOI22_X1 port map( A1 => REGISTERS_21_50_port, A2 => n439, B1 => 
                           REGISTERS_23_50_port, B2 => n402, ZN => n5382);
   U3457 : AOI22_X1 port map( A1 => REGISTERS_17_50_port, A2 => n513, B1 => 
                           REGISTERS_19_50_port, B2 => n476, ZN => n5381);
   U3458 : AOI22_X1 port map( A1 => REGISTERS_20_50_port, A2 => n587, B1 => 
                           REGISTERS_22_50_port, B2 => n550, ZN => n5380);
   U3459 : AOI22_X1 port map( A1 => REGISTERS_16_50_port, A2 => n661, B1 => 
                           REGISTERS_18_50_port, B2 => n624, ZN => n5379);
   U3460 : AND4_X1 port map( A1 => n5382, A2 => n5381, A3 => n5380, A4 => n5379
                           , ZN => n5399);
   U3461 : AOI22_X1 port map( A1 => REGISTERS_29_50_port, A2 => n439, B1 => 
                           REGISTERS_31_50_port, B2 => n402, ZN => n5386);
   U3462 : AOI22_X1 port map( A1 => REGISTERS_25_50_port, A2 => n513, B1 => 
                           REGISTERS_27_50_port, B2 => n476, ZN => n5385);
   U3463 : AOI22_X1 port map( A1 => REGISTERS_28_50_port, A2 => n587, B1 => 
                           REGISTERS_30_50_port, B2 => n550, ZN => n5384);
   U3464 : AOI22_X1 port map( A1 => REGISTERS_24_50_port, A2 => n661, B1 => 
                           REGISTERS_26_50_port, B2 => n624, ZN => n5383);
   U3465 : AND4_X1 port map( A1 => n5386, A2 => n5385, A3 => n5384, A4 => n5383
                           , ZN => n5398);
   U3466 : AOI22_X1 port map( A1 => REGISTERS_5_50_port, A2 => n439, B1 => 
                           REGISTERS_7_50_port, B2 => n402, ZN => n5390);
   U3467 : AOI22_X1 port map( A1 => REGISTERS_1_50_port, A2 => n513, B1 => 
                           REGISTERS_3_50_port, B2 => n476, ZN => n5389);
   U3468 : AOI22_X1 port map( A1 => REGISTERS_4_50_port, A2 => n587, B1 => 
                           REGISTERS_6_50_port, B2 => n550, ZN => n5388);
   U3469 : AOI22_X1 port map( A1 => REGISTERS_0_50_port, A2 => n661, B1 => 
                           REGISTERS_2_50_port, B2 => n624, ZN => n5387);
   U3470 : NAND4_X1 port map( A1 => n5390, A2 => n5389, A3 => n5388, A4 => 
                           n5387, ZN => n5396);
   U3471 : AOI22_X1 port map( A1 => REGISTERS_13_50_port, A2 => n439, B1 => 
                           REGISTERS_15_50_port, B2 => n402, ZN => n5394);
   U3472 : AOI22_X1 port map( A1 => REGISTERS_9_50_port, A2 => n513, B1 => 
                           REGISTERS_11_50_port, B2 => n476, ZN => n5393);
   U3473 : AOI22_X1 port map( A1 => REGISTERS_12_50_port, A2 => n587, B1 => 
                           REGISTERS_14_50_port, B2 => n550, ZN => n5392);
   U3474 : AOI22_X1 port map( A1 => REGISTERS_8_50_port, A2 => n661, B1 => 
                           REGISTERS_10_50_port, B2 => n624, ZN => n5391);
   U3475 : NAND4_X1 port map( A1 => n5394, A2 => n5393, A3 => n5392, A4 => 
                           n5391, ZN => n5395);
   U3476 : AOI22_X1 port map( A1 => n5396, A2 => n23, B1 => n5395, B2 => n22, 
                           ZN => n5397);
   U3477 : OAI221_X1 port map( B1 => n5673, B2 => n5399, C1 => n5671, C2 => 
                           n5398, A => n5397, ZN => N238);
   U3478 : AOI22_X1 port map( A1 => REGISTERS_21_51_port, A2 => n440, B1 => 
                           REGISTERS_23_51_port, B2 => n403, ZN => n5403);
   U3479 : AOI22_X1 port map( A1 => REGISTERS_17_51_port, A2 => n514, B1 => 
                           REGISTERS_19_51_port, B2 => n477, ZN => n5402);
   U3480 : AOI22_X1 port map( A1 => REGISTERS_20_51_port, A2 => n588, B1 => 
                           REGISTERS_22_51_port, B2 => n551, ZN => n5401);
   U3481 : AOI22_X1 port map( A1 => REGISTERS_16_51_port, A2 => n662, B1 => 
                           REGISTERS_18_51_port, B2 => n625, ZN => n5400);
   U3482 : AND4_X1 port map( A1 => n5403, A2 => n5402, A3 => n5401, A4 => n5400
                           , ZN => n5420);
   U3483 : AOI22_X1 port map( A1 => REGISTERS_29_51_port, A2 => n440, B1 => 
                           REGISTERS_31_51_port, B2 => n403, ZN => n5407);
   U3484 : AOI22_X1 port map( A1 => REGISTERS_25_51_port, A2 => n514, B1 => 
                           REGISTERS_27_51_port, B2 => n477, ZN => n5406);
   U3485 : AOI22_X1 port map( A1 => REGISTERS_28_51_port, A2 => n588, B1 => 
                           REGISTERS_30_51_port, B2 => n551, ZN => n5405);
   U3486 : AOI22_X1 port map( A1 => REGISTERS_24_51_port, A2 => n662, B1 => 
                           REGISTERS_26_51_port, B2 => n625, ZN => n5404);
   U3487 : AND4_X1 port map( A1 => n5407, A2 => n5406, A3 => n5405, A4 => n5404
                           , ZN => n5419);
   U3488 : AOI22_X1 port map( A1 => REGISTERS_5_51_port, A2 => n440, B1 => 
                           REGISTERS_7_51_port, B2 => n403, ZN => n5411);
   U3489 : AOI22_X1 port map( A1 => REGISTERS_1_51_port, A2 => n514, B1 => 
                           REGISTERS_3_51_port, B2 => n477, ZN => n5410);
   U3490 : AOI22_X1 port map( A1 => REGISTERS_4_51_port, A2 => n588, B1 => 
                           REGISTERS_6_51_port, B2 => n551, ZN => n5409);
   U3491 : AOI22_X1 port map( A1 => REGISTERS_0_51_port, A2 => n662, B1 => 
                           REGISTERS_2_51_port, B2 => n625, ZN => n5408);
   U3492 : NAND4_X1 port map( A1 => n5411, A2 => n5410, A3 => n5409, A4 => 
                           n5408, ZN => n5417);
   U3493 : AOI22_X1 port map( A1 => REGISTERS_13_51_port, A2 => n440, B1 => 
                           REGISTERS_15_51_port, B2 => n403, ZN => n5415);
   U3494 : AOI22_X1 port map( A1 => REGISTERS_9_51_port, A2 => n514, B1 => 
                           REGISTERS_11_51_port, B2 => n477, ZN => n5414);
   U3495 : AOI22_X1 port map( A1 => REGISTERS_12_51_port, A2 => n588, B1 => 
                           REGISTERS_14_51_port, B2 => n551, ZN => n5413);
   U3496 : AOI22_X1 port map( A1 => REGISTERS_8_51_port, A2 => n662, B1 => 
                           REGISTERS_10_51_port, B2 => n625, ZN => n5412);
   U3497 : NAND4_X1 port map( A1 => n5415, A2 => n5414, A3 => n5413, A4 => 
                           n5412, ZN => n5416);
   U3498 : AOI22_X1 port map( A1 => n5417, A2 => n23, B1 => n5416, B2 => n22, 
                           ZN => n5418);
   U3499 : OAI221_X1 port map( B1 => n5673, B2 => n5420, C1 => n5671, C2 => 
                           n5419, A => n5418, ZN => N237);
   U3500 : AOI22_X1 port map( A1 => REGISTERS_21_52_port, A2 => n440, B1 => 
                           REGISTERS_23_52_port, B2 => n403, ZN => n5424);
   U3501 : AOI22_X1 port map( A1 => REGISTERS_17_52_port, A2 => n514, B1 => 
                           REGISTERS_19_52_port, B2 => n477, ZN => n5423);
   U3502 : AOI22_X1 port map( A1 => REGISTERS_20_52_port, A2 => n588, B1 => 
                           REGISTERS_22_52_port, B2 => n551, ZN => n5422);
   U3503 : AOI22_X1 port map( A1 => REGISTERS_16_52_port, A2 => n662, B1 => 
                           REGISTERS_18_52_port, B2 => n625, ZN => n5421);
   U3504 : AND4_X1 port map( A1 => n5424, A2 => n5423, A3 => n5422, A4 => n5421
                           , ZN => n5441);
   U3505 : AOI22_X1 port map( A1 => REGISTERS_29_52_port, A2 => n440, B1 => 
                           REGISTERS_31_52_port, B2 => n403, ZN => n5428);
   U3506 : AOI22_X1 port map( A1 => REGISTERS_25_52_port, A2 => n514, B1 => 
                           REGISTERS_27_52_port, B2 => n477, ZN => n5427);
   U3507 : AOI22_X1 port map( A1 => REGISTERS_28_52_port, A2 => n588, B1 => 
                           REGISTERS_30_52_port, B2 => n551, ZN => n5426);
   U3508 : AOI22_X1 port map( A1 => REGISTERS_24_52_port, A2 => n662, B1 => 
                           REGISTERS_26_52_port, B2 => n625, ZN => n5425);
   U3509 : AND4_X1 port map( A1 => n5428, A2 => n5427, A3 => n5426, A4 => n5425
                           , ZN => n5440);
   U3510 : AOI22_X1 port map( A1 => REGISTERS_5_52_port, A2 => n440, B1 => 
                           REGISTERS_7_52_port, B2 => n403, ZN => n5432);
   U3511 : AOI22_X1 port map( A1 => REGISTERS_1_52_port, A2 => n514, B1 => 
                           REGISTERS_3_52_port, B2 => n477, ZN => n5431);
   U3512 : AOI22_X1 port map( A1 => REGISTERS_4_52_port, A2 => n588, B1 => 
                           REGISTERS_6_52_port, B2 => n551, ZN => n5430);
   U3513 : AOI22_X1 port map( A1 => REGISTERS_0_52_port, A2 => n662, B1 => 
                           REGISTERS_2_52_port, B2 => n625, ZN => n5429);
   U3514 : NAND4_X1 port map( A1 => n5432, A2 => n5431, A3 => n5430, A4 => 
                           n5429, ZN => n5438);
   U3515 : AOI22_X1 port map( A1 => REGISTERS_13_52_port, A2 => n440, B1 => 
                           REGISTERS_15_52_port, B2 => n403, ZN => n5436);
   U3516 : AOI22_X1 port map( A1 => REGISTERS_9_52_port, A2 => n514, B1 => 
                           REGISTERS_11_52_port, B2 => n477, ZN => n5435);
   U3517 : AOI22_X1 port map( A1 => REGISTERS_12_52_port, A2 => n588, B1 => 
                           REGISTERS_14_52_port, B2 => n551, ZN => n5434);
   U3518 : AOI22_X1 port map( A1 => REGISTERS_8_52_port, A2 => n662, B1 => 
                           REGISTERS_10_52_port, B2 => n625, ZN => n5433);
   U3519 : NAND4_X1 port map( A1 => n5436, A2 => n5435, A3 => n5434, A4 => 
                           n5433, ZN => n5437);
   U3520 : AOI22_X1 port map( A1 => n5438, A2 => n23, B1 => n5437, B2 => n22, 
                           ZN => n5439);
   U3521 : OAI221_X1 port map( B1 => n5673, B2 => n5441, C1 => n5671, C2 => 
                           n5440, A => n5439, ZN => N236);
   U3522 : AOI22_X1 port map( A1 => REGISTERS_21_53_port, A2 => n440, B1 => 
                           REGISTERS_23_53_port, B2 => n403, ZN => n5445);
   U3523 : AOI22_X1 port map( A1 => REGISTERS_17_53_port, A2 => n514, B1 => 
                           REGISTERS_19_53_port, B2 => n477, ZN => n5444);
   U3524 : AOI22_X1 port map( A1 => REGISTERS_20_53_port, A2 => n588, B1 => 
                           REGISTERS_22_53_port, B2 => n551, ZN => n5443);
   U3525 : AOI22_X1 port map( A1 => REGISTERS_16_53_port, A2 => n662, B1 => 
                           REGISTERS_18_53_port, B2 => n625, ZN => n5442);
   U3526 : AND4_X1 port map( A1 => n5445, A2 => n5444, A3 => n5443, A4 => n5442
                           , ZN => n5462);
   U3527 : AOI22_X1 port map( A1 => REGISTERS_29_53_port, A2 => n440, B1 => 
                           REGISTERS_31_53_port, B2 => n403, ZN => n5449);
   U3528 : AOI22_X1 port map( A1 => REGISTERS_25_53_port, A2 => n514, B1 => 
                           REGISTERS_27_53_port, B2 => n477, ZN => n5448);
   U3529 : AOI22_X1 port map( A1 => REGISTERS_28_53_port, A2 => n588, B1 => 
                           REGISTERS_30_53_port, B2 => n551, ZN => n5447);
   U3530 : AOI22_X1 port map( A1 => REGISTERS_24_53_port, A2 => n662, B1 => 
                           REGISTERS_26_53_port, B2 => n625, ZN => n5446);
   U3531 : AND4_X1 port map( A1 => n5449, A2 => n5448, A3 => n5447, A4 => n5446
                           , ZN => n5461);
   U3532 : AOI22_X1 port map( A1 => REGISTERS_5_53_port, A2 => n440, B1 => 
                           REGISTERS_7_53_port, B2 => n403, ZN => n5453);
   U3533 : AOI22_X1 port map( A1 => REGISTERS_1_53_port, A2 => n514, B1 => 
                           REGISTERS_3_53_port, B2 => n477, ZN => n5452);
   U3534 : AOI22_X1 port map( A1 => REGISTERS_4_53_port, A2 => n588, B1 => 
                           REGISTERS_6_53_port, B2 => n551, ZN => n5451);
   U3535 : AOI22_X1 port map( A1 => REGISTERS_0_53_port, A2 => n662, B1 => 
                           REGISTERS_2_53_port, B2 => n625, ZN => n5450);
   U3536 : NAND4_X1 port map( A1 => n5453, A2 => n5452, A3 => n5451, A4 => 
                           n5450, ZN => n5459);
   U3537 : AOI22_X1 port map( A1 => REGISTERS_13_53_port, A2 => n440, B1 => 
                           REGISTERS_15_53_port, B2 => n403, ZN => n5457);
   U3538 : AOI22_X1 port map( A1 => REGISTERS_9_53_port, A2 => n514, B1 => 
                           REGISTERS_11_53_port, B2 => n477, ZN => n5456);
   U3539 : AOI22_X1 port map( A1 => REGISTERS_12_53_port, A2 => n588, B1 => 
                           REGISTERS_14_53_port, B2 => n551, ZN => n5455);
   U3540 : AOI22_X1 port map( A1 => REGISTERS_8_53_port, A2 => n662, B1 => 
                           REGISTERS_10_53_port, B2 => n625, ZN => n5454);
   U3541 : NAND4_X1 port map( A1 => n5457, A2 => n5456, A3 => n5455, A4 => 
                           n5454, ZN => n5458);
   U3542 : AOI22_X1 port map( A1 => n5459, A2 => n23, B1 => n5458, B2 => n22, 
                           ZN => n5460);
   U3543 : OAI221_X1 port map( B1 => n5673, B2 => n5462, C1 => n5671, C2 => 
                           n5461, A => n5460, ZN => N235);
   U3544 : AOI22_X1 port map( A1 => REGISTERS_21_54_port, A2 => n441, B1 => 
                           REGISTERS_23_54_port, B2 => n404, ZN => n5466);
   U3545 : AOI22_X1 port map( A1 => REGISTERS_17_54_port, A2 => n515, B1 => 
                           REGISTERS_19_54_port, B2 => n478, ZN => n5465);
   U3546 : AOI22_X1 port map( A1 => REGISTERS_20_54_port, A2 => n589, B1 => 
                           REGISTERS_22_54_port, B2 => n552, ZN => n5464);
   U3547 : AOI22_X1 port map( A1 => REGISTERS_16_54_port, A2 => n663, B1 => 
                           REGISTERS_18_54_port, B2 => n626, ZN => n5463);
   U3548 : AND4_X1 port map( A1 => n5466, A2 => n5465, A3 => n5464, A4 => n5463
                           , ZN => n5483);
   U3549 : AOI22_X1 port map( A1 => REGISTERS_29_54_port, A2 => n441, B1 => 
                           REGISTERS_31_54_port, B2 => n404, ZN => n5470);
   U3550 : AOI22_X1 port map( A1 => REGISTERS_25_54_port, A2 => n515, B1 => 
                           REGISTERS_27_54_port, B2 => n478, ZN => n5469);
   U3551 : AOI22_X1 port map( A1 => REGISTERS_28_54_port, A2 => n589, B1 => 
                           REGISTERS_30_54_port, B2 => n552, ZN => n5468);
   U3552 : AOI22_X1 port map( A1 => REGISTERS_24_54_port, A2 => n663, B1 => 
                           REGISTERS_26_54_port, B2 => n626, ZN => n5467);
   U3553 : AND4_X1 port map( A1 => n5470, A2 => n5469, A3 => n5468, A4 => n5467
                           , ZN => n5482);
   U3554 : AOI22_X1 port map( A1 => REGISTERS_5_54_port, A2 => n441, B1 => 
                           REGISTERS_7_54_port, B2 => n404, ZN => n5474);
   U3555 : AOI22_X1 port map( A1 => REGISTERS_1_54_port, A2 => n515, B1 => 
                           REGISTERS_3_54_port, B2 => n478, ZN => n5473);
   U3556 : AOI22_X1 port map( A1 => REGISTERS_4_54_port, A2 => n589, B1 => 
                           REGISTERS_6_54_port, B2 => n552, ZN => n5472);
   U3557 : AOI22_X1 port map( A1 => REGISTERS_0_54_port, A2 => n663, B1 => 
                           REGISTERS_2_54_port, B2 => n626, ZN => n5471);
   U3558 : NAND4_X1 port map( A1 => n5474, A2 => n5473, A3 => n5472, A4 => 
                           n5471, ZN => n5480);
   U3559 : AOI22_X1 port map( A1 => REGISTERS_13_54_port, A2 => n441, B1 => 
                           REGISTERS_15_54_port, B2 => n404, ZN => n5478);
   U3560 : AOI22_X1 port map( A1 => REGISTERS_9_54_port, A2 => n515, B1 => 
                           REGISTERS_11_54_port, B2 => n478, ZN => n5477);
   U3561 : AOI22_X1 port map( A1 => REGISTERS_12_54_port, A2 => n589, B1 => 
                           REGISTERS_14_54_port, B2 => n552, ZN => n5476);
   U3562 : AOI22_X1 port map( A1 => REGISTERS_8_54_port, A2 => n663, B1 => 
                           REGISTERS_10_54_port, B2 => n626, ZN => n5475);
   U3563 : NAND4_X1 port map( A1 => n5478, A2 => n5477, A3 => n5476, A4 => 
                           n5475, ZN => n5479);
   U3564 : AOI22_X1 port map( A1 => n5480, A2 => n23, B1 => n5479, B2 => n22, 
                           ZN => n5481);
   U3565 : OAI221_X1 port map( B1 => n5673, B2 => n5483, C1 => n5671, C2 => 
                           n5482, A => n5481, ZN => N234);
   U3566 : AOI22_X1 port map( A1 => REGISTERS_21_55_port, A2 => n441, B1 => 
                           REGISTERS_23_55_port, B2 => n404, ZN => n5487);
   U3567 : AOI22_X1 port map( A1 => REGISTERS_17_55_port, A2 => n515, B1 => 
                           REGISTERS_19_55_port, B2 => n478, ZN => n5486);
   U3568 : AOI22_X1 port map( A1 => REGISTERS_20_55_port, A2 => n589, B1 => 
                           REGISTERS_22_55_port, B2 => n552, ZN => n5485);
   U3569 : AOI22_X1 port map( A1 => REGISTERS_16_55_port, A2 => n663, B1 => 
                           REGISTERS_18_55_port, B2 => n626, ZN => n5484);
   U3570 : AND4_X1 port map( A1 => n5487, A2 => n5486, A3 => n5485, A4 => n5484
                           , ZN => n5504);
   U3571 : AOI22_X1 port map( A1 => REGISTERS_29_55_port, A2 => n441, B1 => 
                           REGISTERS_31_55_port, B2 => n404, ZN => n5491);
   U3572 : AOI22_X1 port map( A1 => REGISTERS_25_55_port, A2 => n515, B1 => 
                           REGISTERS_27_55_port, B2 => n478, ZN => n5490);
   U3573 : AOI22_X1 port map( A1 => REGISTERS_28_55_port, A2 => n589, B1 => 
                           REGISTERS_30_55_port, B2 => n552, ZN => n5489);
   U3574 : AOI22_X1 port map( A1 => REGISTERS_24_55_port, A2 => n663, B1 => 
                           REGISTERS_26_55_port, B2 => n626, ZN => n5488);
   U3575 : AND4_X1 port map( A1 => n5491, A2 => n5490, A3 => n5489, A4 => n5488
                           , ZN => n5503);
   U3576 : AOI22_X1 port map( A1 => REGISTERS_5_55_port, A2 => n441, B1 => 
                           REGISTERS_7_55_port, B2 => n404, ZN => n5495);
   U3577 : AOI22_X1 port map( A1 => REGISTERS_1_55_port, A2 => n515, B1 => 
                           REGISTERS_3_55_port, B2 => n478, ZN => n5494);
   U3578 : AOI22_X1 port map( A1 => REGISTERS_4_55_port, A2 => n589, B1 => 
                           REGISTERS_6_55_port, B2 => n552, ZN => n5493);
   U3579 : AOI22_X1 port map( A1 => REGISTERS_0_55_port, A2 => n663, B1 => 
                           REGISTERS_2_55_port, B2 => n626, ZN => n5492);
   U3580 : NAND4_X1 port map( A1 => n5495, A2 => n5494, A3 => n5493, A4 => 
                           n5492, ZN => n5501);
   U3581 : AOI22_X1 port map( A1 => REGISTERS_13_55_port, A2 => n441, B1 => 
                           REGISTERS_15_55_port, B2 => n404, ZN => n5499);
   U3582 : AOI22_X1 port map( A1 => REGISTERS_9_55_port, A2 => n515, B1 => 
                           REGISTERS_11_55_port, B2 => n478, ZN => n5498);
   U3583 : AOI22_X1 port map( A1 => REGISTERS_12_55_port, A2 => n589, B1 => 
                           REGISTERS_14_55_port, B2 => n552, ZN => n5497);
   U3584 : AOI22_X1 port map( A1 => REGISTERS_8_55_port, A2 => n663, B1 => 
                           REGISTERS_10_55_port, B2 => n626, ZN => n5496);
   U3585 : NAND4_X1 port map( A1 => n5499, A2 => n5498, A3 => n5497, A4 => 
                           n5496, ZN => n5500);
   U3586 : AOI22_X1 port map( A1 => n5501, A2 => n23, B1 => n5500, B2 => n22, 
                           ZN => n5502);
   U3587 : OAI221_X1 port map( B1 => n5673, B2 => n5504, C1 => n5671, C2 => 
                           n5503, A => n5502, ZN => N233);
   U3588 : AOI22_X1 port map( A1 => REGISTERS_21_56_port, A2 => n441, B1 => 
                           REGISTERS_23_56_port, B2 => n404, ZN => n5508);
   U3589 : AOI22_X1 port map( A1 => REGISTERS_17_56_port, A2 => n515, B1 => 
                           REGISTERS_19_56_port, B2 => n478, ZN => n5507);
   U3590 : AOI22_X1 port map( A1 => REGISTERS_20_56_port, A2 => n589, B1 => 
                           REGISTERS_22_56_port, B2 => n552, ZN => n5506);
   U3591 : AOI22_X1 port map( A1 => REGISTERS_16_56_port, A2 => n663, B1 => 
                           REGISTERS_18_56_port, B2 => n626, ZN => n5505);
   U3592 : AND4_X1 port map( A1 => n5508, A2 => n5507, A3 => n5506, A4 => n5505
                           , ZN => n5525);
   U3593 : AOI22_X1 port map( A1 => REGISTERS_29_56_port, A2 => n441, B1 => 
                           REGISTERS_31_56_port, B2 => n404, ZN => n5512);
   U3594 : AOI22_X1 port map( A1 => REGISTERS_25_56_port, A2 => n515, B1 => 
                           REGISTERS_27_56_port, B2 => n478, ZN => n5511);
   U3595 : AOI22_X1 port map( A1 => REGISTERS_28_56_port, A2 => n589, B1 => 
                           REGISTERS_30_56_port, B2 => n552, ZN => n5510);
   U3596 : AOI22_X1 port map( A1 => REGISTERS_24_56_port, A2 => n663, B1 => 
                           REGISTERS_26_56_port, B2 => n626, ZN => n5509);
   U3597 : AND4_X1 port map( A1 => n5512, A2 => n5511, A3 => n5510, A4 => n5509
                           , ZN => n5524);
   U3598 : AOI22_X1 port map( A1 => REGISTERS_5_56_port, A2 => n441, B1 => 
                           REGISTERS_7_56_port, B2 => n404, ZN => n5516);
   U3599 : AOI22_X1 port map( A1 => REGISTERS_1_56_port, A2 => n515, B1 => 
                           REGISTERS_3_56_port, B2 => n478, ZN => n5515);
   U3600 : AOI22_X1 port map( A1 => REGISTERS_4_56_port, A2 => n589, B1 => 
                           REGISTERS_6_56_port, B2 => n552, ZN => n5514);
   U3601 : AOI22_X1 port map( A1 => REGISTERS_0_56_port, A2 => n663, B1 => 
                           REGISTERS_2_56_port, B2 => n626, ZN => n5513);
   U3602 : NAND4_X1 port map( A1 => n5516, A2 => n5515, A3 => n5514, A4 => 
                           n5513, ZN => n5522);
   U3603 : AOI22_X1 port map( A1 => REGISTERS_13_56_port, A2 => n441, B1 => 
                           REGISTERS_15_56_port, B2 => n404, ZN => n5520);
   U3604 : AOI22_X1 port map( A1 => REGISTERS_9_56_port, A2 => n515, B1 => 
                           REGISTERS_11_56_port, B2 => n478, ZN => n5519);
   U3605 : AOI22_X1 port map( A1 => REGISTERS_12_56_port, A2 => n589, B1 => 
                           REGISTERS_14_56_port, B2 => n552, ZN => n5518);
   U3606 : AOI22_X1 port map( A1 => REGISTERS_8_56_port, A2 => n663, B1 => 
                           REGISTERS_10_56_port, B2 => n626, ZN => n5517);
   U3607 : NAND4_X1 port map( A1 => n5520, A2 => n5519, A3 => n5518, A4 => 
                           n5517, ZN => n5521);
   U3608 : AOI22_X1 port map( A1 => n5522, A2 => n23, B1 => n5521, B2 => n22, 
                           ZN => n5523);
   U3609 : OAI221_X1 port map( B1 => n5673, B2 => n5525, C1 => n5671, C2 => 
                           n5524, A => n5523, ZN => N232);
   U3610 : AOI22_X1 port map( A1 => REGISTERS_21_57_port, A2 => n442, B1 => 
                           REGISTERS_23_57_port, B2 => n405, ZN => n5529);
   U3611 : AOI22_X1 port map( A1 => REGISTERS_17_57_port, A2 => n516, B1 => 
                           REGISTERS_19_57_port, B2 => n479, ZN => n5528);
   U3612 : AOI22_X1 port map( A1 => REGISTERS_20_57_port, A2 => n590, B1 => 
                           REGISTERS_22_57_port, B2 => n553, ZN => n5527);
   U3613 : AOI22_X1 port map( A1 => REGISTERS_16_57_port, A2 => n664, B1 => 
                           REGISTERS_18_57_port, B2 => n627, ZN => n5526);
   U3614 : AND4_X1 port map( A1 => n5529, A2 => n5528, A3 => n5527, A4 => n5526
                           , ZN => n5546);
   U3615 : AOI22_X1 port map( A1 => REGISTERS_29_57_port, A2 => n442, B1 => 
                           REGISTERS_31_57_port, B2 => n405, ZN => n5533);
   U3616 : AOI22_X1 port map( A1 => REGISTERS_25_57_port, A2 => n516, B1 => 
                           REGISTERS_27_57_port, B2 => n479, ZN => n5532);
   U3617 : AOI22_X1 port map( A1 => REGISTERS_28_57_port, A2 => n590, B1 => 
                           REGISTERS_30_57_port, B2 => n553, ZN => n5531);
   U3618 : AOI22_X1 port map( A1 => REGISTERS_24_57_port, A2 => n664, B1 => 
                           REGISTERS_26_57_port, B2 => n627, ZN => n5530);
   U3619 : AND4_X1 port map( A1 => n5533, A2 => n5532, A3 => n5531, A4 => n5530
                           , ZN => n5545);
   U3620 : AOI22_X1 port map( A1 => REGISTERS_5_57_port, A2 => n442, B1 => 
                           REGISTERS_7_57_port, B2 => n405, ZN => n5537);
   U3621 : AOI22_X1 port map( A1 => REGISTERS_1_57_port, A2 => n516, B1 => 
                           REGISTERS_3_57_port, B2 => n479, ZN => n5536);
   U3622 : AOI22_X1 port map( A1 => REGISTERS_4_57_port, A2 => n590, B1 => 
                           REGISTERS_6_57_port, B2 => n553, ZN => n5535);
   U3623 : AOI22_X1 port map( A1 => REGISTERS_0_57_port, A2 => n664, B1 => 
                           REGISTERS_2_57_port, B2 => n627, ZN => n5534);
   U3624 : NAND4_X1 port map( A1 => n5537, A2 => n5536, A3 => n5535, A4 => 
                           n5534, ZN => n5543);
   U3625 : AOI22_X1 port map( A1 => REGISTERS_13_57_port, A2 => n442, B1 => 
                           REGISTERS_15_57_port, B2 => n405, ZN => n5541);
   U3626 : AOI22_X1 port map( A1 => REGISTERS_9_57_port, A2 => n516, B1 => 
                           REGISTERS_11_57_port, B2 => n479, ZN => n5540);
   U3627 : AOI22_X1 port map( A1 => REGISTERS_12_57_port, A2 => n590, B1 => 
                           REGISTERS_14_57_port, B2 => n553, ZN => n5539);
   U3628 : AOI22_X1 port map( A1 => REGISTERS_8_57_port, A2 => n664, B1 => 
                           REGISTERS_10_57_port, B2 => n627, ZN => n5538);
   U3629 : NAND4_X1 port map( A1 => n5541, A2 => n5540, A3 => n5539, A4 => 
                           n5538, ZN => n5542);
   U3630 : AOI22_X1 port map( A1 => n5543, A2 => n23, B1 => n5542, B2 => n22, 
                           ZN => n5544);
   U3631 : OAI221_X1 port map( B1 => n5673, B2 => n5546, C1 => n5671, C2 => 
                           n5545, A => n5544, ZN => N231);
   U3632 : AOI22_X1 port map( A1 => REGISTERS_21_58_port, A2 => n442, B1 => 
                           REGISTERS_23_58_port, B2 => n405, ZN => n5550);
   U3633 : AOI22_X1 port map( A1 => REGISTERS_17_58_port, A2 => n516, B1 => 
                           REGISTERS_19_58_port, B2 => n479, ZN => n5549);
   U3634 : AOI22_X1 port map( A1 => REGISTERS_20_58_port, A2 => n590, B1 => 
                           REGISTERS_22_58_port, B2 => n553, ZN => n5548);
   U3635 : AOI22_X1 port map( A1 => REGISTERS_16_58_port, A2 => n664, B1 => 
                           REGISTERS_18_58_port, B2 => n627, ZN => n5547);
   U3636 : AND4_X1 port map( A1 => n5550, A2 => n5549, A3 => n5548, A4 => n5547
                           , ZN => n5567);
   U3637 : AOI22_X1 port map( A1 => REGISTERS_29_58_port, A2 => n442, B1 => 
                           REGISTERS_31_58_port, B2 => n405, ZN => n5554);
   U3638 : AOI22_X1 port map( A1 => REGISTERS_25_58_port, A2 => n516, B1 => 
                           REGISTERS_27_58_port, B2 => n479, ZN => n5553);
   U3639 : AOI22_X1 port map( A1 => REGISTERS_28_58_port, A2 => n590, B1 => 
                           REGISTERS_30_58_port, B2 => n553, ZN => n5552);
   U3640 : AOI22_X1 port map( A1 => REGISTERS_24_58_port, A2 => n664, B1 => 
                           REGISTERS_26_58_port, B2 => n627, ZN => n5551);
   U3641 : AND4_X1 port map( A1 => n5554, A2 => n5553, A3 => n5552, A4 => n5551
                           , ZN => n5566);
   U3642 : AOI22_X1 port map( A1 => REGISTERS_5_58_port, A2 => n442, B1 => 
                           REGISTERS_7_58_port, B2 => n405, ZN => n5558);
   U3643 : AOI22_X1 port map( A1 => REGISTERS_1_58_port, A2 => n516, B1 => 
                           REGISTERS_3_58_port, B2 => n479, ZN => n5557);
   U3644 : AOI22_X1 port map( A1 => REGISTERS_4_58_port, A2 => n590, B1 => 
                           REGISTERS_6_58_port, B2 => n553, ZN => n5556);
   U3645 : AOI22_X1 port map( A1 => REGISTERS_0_58_port, A2 => n664, B1 => 
                           REGISTERS_2_58_port, B2 => n627, ZN => n5555);
   U3646 : NAND4_X1 port map( A1 => n5558, A2 => n5557, A3 => n5556, A4 => 
                           n5555, ZN => n5564);
   U3647 : AOI22_X1 port map( A1 => REGISTERS_13_58_port, A2 => n442, B1 => 
                           REGISTERS_15_58_port, B2 => n405, ZN => n5562);
   U3648 : AOI22_X1 port map( A1 => REGISTERS_9_58_port, A2 => n516, B1 => 
                           REGISTERS_11_58_port, B2 => n479, ZN => n5561);
   U3649 : AOI22_X1 port map( A1 => REGISTERS_12_58_port, A2 => n590, B1 => 
                           REGISTERS_14_58_port, B2 => n553, ZN => n5560);
   U3650 : AOI22_X1 port map( A1 => REGISTERS_8_58_port, A2 => n664, B1 => 
                           REGISTERS_10_58_port, B2 => n627, ZN => n5559);
   U3651 : NAND4_X1 port map( A1 => n5562, A2 => n5561, A3 => n5560, A4 => 
                           n5559, ZN => n5563);
   U3652 : AOI22_X1 port map( A1 => n5564, A2 => n23, B1 => n5563, B2 => n22, 
                           ZN => n5565);
   U3653 : OAI221_X1 port map( B1 => n5673, B2 => n5567, C1 => n5671, C2 => 
                           n5566, A => n5565, ZN => N230);
   U3654 : AOI22_X1 port map( A1 => REGISTERS_21_59_port, A2 => n442, B1 => 
                           REGISTERS_23_59_port, B2 => n405, ZN => n5571);
   U3655 : AOI22_X1 port map( A1 => REGISTERS_17_59_port, A2 => n516, B1 => 
                           REGISTERS_19_59_port, B2 => n479, ZN => n5570);
   U3656 : AOI22_X1 port map( A1 => REGISTERS_20_59_port, A2 => n590, B1 => 
                           REGISTERS_22_59_port, B2 => n553, ZN => n5569);
   U3657 : AOI22_X1 port map( A1 => REGISTERS_16_59_port, A2 => n664, B1 => 
                           REGISTERS_18_59_port, B2 => n627, ZN => n5568);
   U3658 : AND4_X1 port map( A1 => n5571, A2 => n5570, A3 => n5569, A4 => n5568
                           , ZN => n5588);
   U3659 : AOI22_X1 port map( A1 => REGISTERS_29_59_port, A2 => n442, B1 => 
                           REGISTERS_31_59_port, B2 => n405, ZN => n5575);
   U3660 : AOI22_X1 port map( A1 => REGISTERS_25_59_port, A2 => n516, B1 => 
                           REGISTERS_27_59_port, B2 => n479, ZN => n5574);
   U3661 : AOI22_X1 port map( A1 => REGISTERS_28_59_port, A2 => n590, B1 => 
                           REGISTERS_30_59_port, B2 => n553, ZN => n5573);
   U3662 : AOI22_X1 port map( A1 => REGISTERS_24_59_port, A2 => n664, B1 => 
                           REGISTERS_26_59_port, B2 => n627, ZN => n5572);
   U3663 : AND4_X1 port map( A1 => n5575, A2 => n5574, A3 => n5573, A4 => n5572
                           , ZN => n5587);
   U3664 : AOI22_X1 port map( A1 => REGISTERS_5_59_port, A2 => n442, B1 => 
                           REGISTERS_7_59_port, B2 => n405, ZN => n5579);
   U3665 : AOI22_X1 port map( A1 => REGISTERS_1_59_port, A2 => n516, B1 => 
                           REGISTERS_3_59_port, B2 => n479, ZN => n5578);
   U3666 : AOI22_X1 port map( A1 => REGISTERS_4_59_port, A2 => n590, B1 => 
                           REGISTERS_6_59_port, B2 => n553, ZN => n5577);
   U3667 : AOI22_X1 port map( A1 => REGISTERS_0_59_port, A2 => n664, B1 => 
                           REGISTERS_2_59_port, B2 => n627, ZN => n5576);
   U3668 : NAND4_X1 port map( A1 => n5579, A2 => n5578, A3 => n5577, A4 => 
                           n5576, ZN => n5585);
   U3669 : AOI22_X1 port map( A1 => REGISTERS_13_59_port, A2 => n442, B1 => 
                           REGISTERS_15_59_port, B2 => n405, ZN => n5583);
   U3670 : AOI22_X1 port map( A1 => REGISTERS_9_59_port, A2 => n516, B1 => 
                           REGISTERS_11_59_port, B2 => n479, ZN => n5582);
   U3671 : AOI22_X1 port map( A1 => REGISTERS_12_59_port, A2 => n590, B1 => 
                           REGISTERS_14_59_port, B2 => n553, ZN => n5581);
   U3672 : AOI22_X1 port map( A1 => REGISTERS_8_59_port, A2 => n664, B1 => 
                           REGISTERS_10_59_port, B2 => n627, ZN => n5580);
   U3673 : NAND4_X1 port map( A1 => n5583, A2 => n5582, A3 => n5581, A4 => 
                           n5580, ZN => n5584);
   U3674 : AOI22_X1 port map( A1 => n5585, A2 => n23, B1 => n5584, B2 => n22, 
                           ZN => n5586);
   U3675 : OAI221_X1 port map( B1 => n5673, B2 => n5588, C1 => n5671, C2 => 
                           n5587, A => n5586, ZN => N229);
   U3676 : AOI22_X1 port map( A1 => REGISTERS_21_60_port, A2 => n443, B1 => 
                           REGISTERS_23_60_port, B2 => n406, ZN => n5592);
   U3677 : AOI22_X1 port map( A1 => REGISTERS_17_60_port, A2 => n517, B1 => 
                           REGISTERS_19_60_port, B2 => n480, ZN => n5591);
   U3678 : AOI22_X1 port map( A1 => REGISTERS_20_60_port, A2 => n591, B1 => 
                           REGISTERS_22_60_port, B2 => n554, ZN => n5590);
   U3679 : AOI22_X1 port map( A1 => REGISTERS_16_60_port, A2 => n665, B1 => 
                           REGISTERS_18_60_port, B2 => n628, ZN => n5589);
   U3680 : AND4_X1 port map( A1 => n5592, A2 => n5591, A3 => n5590, A4 => n5589
                           , ZN => n5609);
   U3681 : AOI22_X1 port map( A1 => REGISTERS_29_60_port, A2 => n443, B1 => 
                           REGISTERS_31_60_port, B2 => n406, ZN => n5596);
   U3682 : AOI22_X1 port map( A1 => REGISTERS_25_60_port, A2 => n517, B1 => 
                           REGISTERS_27_60_port, B2 => n480, ZN => n5595);
   U3683 : AOI22_X1 port map( A1 => REGISTERS_28_60_port, A2 => n591, B1 => 
                           REGISTERS_30_60_port, B2 => n554, ZN => n5594);
   U3684 : AOI22_X1 port map( A1 => REGISTERS_24_60_port, A2 => n665, B1 => 
                           REGISTERS_26_60_port, B2 => n628, ZN => n5593);
   U3685 : AND4_X1 port map( A1 => n5596, A2 => n5595, A3 => n5594, A4 => n5593
                           , ZN => n5608);
   U3686 : AOI22_X1 port map( A1 => REGISTERS_5_60_port, A2 => n443, B1 => 
                           REGISTERS_7_60_port, B2 => n406, ZN => n5600);
   U3687 : AOI22_X1 port map( A1 => REGISTERS_1_60_port, A2 => n517, B1 => 
                           REGISTERS_3_60_port, B2 => n480, ZN => n5599);
   U3688 : AOI22_X1 port map( A1 => REGISTERS_4_60_port, A2 => n591, B1 => 
                           REGISTERS_6_60_port, B2 => n554, ZN => n5598);
   U3689 : AOI22_X1 port map( A1 => REGISTERS_0_60_port, A2 => n665, B1 => 
                           REGISTERS_2_60_port, B2 => n628, ZN => n5597);
   U3690 : NAND4_X1 port map( A1 => n5600, A2 => n5599, A3 => n5598, A4 => 
                           n5597, ZN => n5606);
   U3691 : AOI22_X1 port map( A1 => REGISTERS_13_60_port, A2 => n443, B1 => 
                           REGISTERS_15_60_port, B2 => n406, ZN => n5604);
   U3692 : AOI22_X1 port map( A1 => REGISTERS_9_60_port, A2 => n517, B1 => 
                           REGISTERS_11_60_port, B2 => n480, ZN => n5603);
   U3693 : AOI22_X1 port map( A1 => REGISTERS_12_60_port, A2 => n591, B1 => 
                           REGISTERS_14_60_port, B2 => n554, ZN => n5602);
   U3694 : AOI22_X1 port map( A1 => REGISTERS_8_60_port, A2 => n665, B1 => 
                           REGISTERS_10_60_port, B2 => n628, ZN => n5601);
   U3695 : NAND4_X1 port map( A1 => n5604, A2 => n5603, A3 => n5602, A4 => 
                           n5601, ZN => n5605);
   U3696 : AOI22_X1 port map( A1 => n5606, A2 => n23, B1 => n5605, B2 => n22, 
                           ZN => n5607);
   U3697 : OAI221_X1 port map( B1 => n5673, B2 => n5609, C1 => n5671, C2 => 
                           n5608, A => n5607, ZN => N228);
   U3698 : AOI22_X1 port map( A1 => REGISTERS_21_61_port, A2 => n443, B1 => 
                           REGISTERS_23_61_port, B2 => n406, ZN => n5613);
   U3699 : AOI22_X1 port map( A1 => REGISTERS_17_61_port, A2 => n517, B1 => 
                           REGISTERS_19_61_port, B2 => n480, ZN => n5612);
   U3700 : AOI22_X1 port map( A1 => REGISTERS_20_61_port, A2 => n591, B1 => 
                           REGISTERS_22_61_port, B2 => n554, ZN => n5611);
   U3701 : AOI22_X1 port map( A1 => REGISTERS_16_61_port, A2 => n665, B1 => 
                           REGISTERS_18_61_port, B2 => n628, ZN => n5610);
   U3702 : AND4_X1 port map( A1 => n5613, A2 => n5612, A3 => n5611, A4 => n5610
                           , ZN => n5630);
   U3703 : AOI22_X1 port map( A1 => REGISTERS_29_61_port, A2 => n443, B1 => 
                           REGISTERS_31_61_port, B2 => n406, ZN => n5617);
   U3704 : AOI22_X1 port map( A1 => REGISTERS_25_61_port, A2 => n517, B1 => 
                           REGISTERS_27_61_port, B2 => n480, ZN => n5616);
   U3705 : AOI22_X1 port map( A1 => REGISTERS_28_61_port, A2 => n591, B1 => 
                           REGISTERS_30_61_port, B2 => n554, ZN => n5615);
   U3706 : AOI22_X1 port map( A1 => REGISTERS_24_61_port, A2 => n665, B1 => 
                           REGISTERS_26_61_port, B2 => n628, ZN => n5614);
   U3707 : AND4_X1 port map( A1 => n5617, A2 => n5616, A3 => n5615, A4 => n5614
                           , ZN => n5629);
   U3708 : AOI22_X1 port map( A1 => REGISTERS_5_61_port, A2 => n443, B1 => 
                           REGISTERS_7_61_port, B2 => n406, ZN => n5621);
   U3709 : AOI22_X1 port map( A1 => REGISTERS_1_61_port, A2 => n517, B1 => 
                           REGISTERS_3_61_port, B2 => n480, ZN => n5620);
   U3710 : AOI22_X1 port map( A1 => REGISTERS_4_61_port, A2 => n591, B1 => 
                           REGISTERS_6_61_port, B2 => n554, ZN => n5619);
   U3711 : AOI22_X1 port map( A1 => REGISTERS_0_61_port, A2 => n665, B1 => 
                           REGISTERS_2_61_port, B2 => n628, ZN => n5618);
   U3712 : NAND4_X1 port map( A1 => n5621, A2 => n5620, A3 => n5619, A4 => 
                           n5618, ZN => n5627);
   U3713 : AOI22_X1 port map( A1 => REGISTERS_13_61_port, A2 => n443, B1 => 
                           REGISTERS_15_61_port, B2 => n406, ZN => n5625);
   U3714 : AOI22_X1 port map( A1 => REGISTERS_9_61_port, A2 => n517, B1 => 
                           REGISTERS_11_61_port, B2 => n480, ZN => n5624);
   U3715 : AOI22_X1 port map( A1 => REGISTERS_12_61_port, A2 => n591, B1 => 
                           REGISTERS_14_61_port, B2 => n554, ZN => n5623);
   U3716 : AOI22_X1 port map( A1 => REGISTERS_8_61_port, A2 => n665, B1 => 
                           REGISTERS_10_61_port, B2 => n628, ZN => n5622);
   U3717 : NAND4_X1 port map( A1 => n5625, A2 => n5624, A3 => n5623, A4 => 
                           n5622, ZN => n5626);
   U3718 : AOI22_X1 port map( A1 => n5627, A2 => n23, B1 => n5626, B2 => n22, 
                           ZN => n5628);
   U3719 : OAI221_X1 port map( B1 => n5673, B2 => n5630, C1 => n5671, C2 => 
                           n5629, A => n5628, ZN => N227);
   U3720 : AOI22_X1 port map( A1 => REGISTERS_21_62_port, A2 => n443, B1 => 
                           REGISTERS_23_62_port, B2 => n406, ZN => n5634);
   U3721 : AOI22_X1 port map( A1 => REGISTERS_17_62_port, A2 => n517, B1 => 
                           REGISTERS_19_62_port, B2 => n480, ZN => n5633);
   U3722 : AOI22_X1 port map( A1 => REGISTERS_20_62_port, A2 => n591, B1 => 
                           REGISTERS_22_62_port, B2 => n554, ZN => n5632);
   U3723 : AOI22_X1 port map( A1 => REGISTERS_16_62_port, A2 => n665, B1 => 
                           REGISTERS_18_62_port, B2 => n628, ZN => n5631);
   U3724 : AND4_X1 port map( A1 => n5634, A2 => n5633, A3 => n5632, A4 => n5631
                           , ZN => n5651);
   U3725 : AOI22_X1 port map( A1 => REGISTERS_29_62_port, A2 => n443, B1 => 
                           REGISTERS_31_62_port, B2 => n406, ZN => n5638);
   U3726 : AOI22_X1 port map( A1 => REGISTERS_25_62_port, A2 => n517, B1 => 
                           REGISTERS_27_62_port, B2 => n480, ZN => n5637);
   U3727 : AOI22_X1 port map( A1 => REGISTERS_28_62_port, A2 => n591, B1 => 
                           REGISTERS_30_62_port, B2 => n554, ZN => n5636);
   U3728 : AOI22_X1 port map( A1 => REGISTERS_24_62_port, A2 => n665, B1 => 
                           REGISTERS_26_62_port, B2 => n628, ZN => n5635);
   U3729 : AND4_X1 port map( A1 => n5638, A2 => n5637, A3 => n5636, A4 => n5635
                           , ZN => n5650);
   U3730 : AOI22_X1 port map( A1 => REGISTERS_5_62_port, A2 => n443, B1 => 
                           REGISTERS_7_62_port, B2 => n406, ZN => n5642);
   U3731 : AOI22_X1 port map( A1 => REGISTERS_1_62_port, A2 => n517, B1 => 
                           REGISTERS_3_62_port, B2 => n480, ZN => n5641);
   U3732 : AOI22_X1 port map( A1 => REGISTERS_4_62_port, A2 => n591, B1 => 
                           REGISTERS_6_62_port, B2 => n554, ZN => n5640);
   U3733 : AOI22_X1 port map( A1 => REGISTERS_0_62_port, A2 => n665, B1 => 
                           REGISTERS_2_62_port, B2 => n628, ZN => n5639);
   U3734 : NAND4_X1 port map( A1 => n5642, A2 => n5641, A3 => n5640, A4 => 
                           n5639, ZN => n5648);
   U3735 : AOI22_X1 port map( A1 => REGISTERS_13_62_port, A2 => n443, B1 => 
                           REGISTERS_15_62_port, B2 => n406, ZN => n5646);
   U3736 : AOI22_X1 port map( A1 => REGISTERS_9_62_port, A2 => n517, B1 => 
                           REGISTERS_11_62_port, B2 => n480, ZN => n5645);
   U3737 : AOI22_X1 port map( A1 => REGISTERS_12_62_port, A2 => n591, B1 => 
                           REGISTERS_14_62_port, B2 => n554, ZN => n5644);
   U3738 : AOI22_X1 port map( A1 => REGISTERS_8_62_port, A2 => n665, B1 => 
                           REGISTERS_10_62_port, B2 => n628, ZN => n5643);
   U3739 : NAND4_X1 port map( A1 => n5646, A2 => n5645, A3 => n5644, A4 => 
                           n5643, ZN => n5647);
   U3740 : AOI22_X1 port map( A1 => n5648, A2 => n23, B1 => n5647, B2 => n22, 
                           ZN => n5649);
   U3741 : OAI221_X1 port map( B1 => n5673, B2 => n5651, C1 => n5671, C2 => 
                           n5650, A => n5649, ZN => N226);
   U3742 : AOI22_X1 port map( A1 => REGISTERS_21_63_port, A2 => n444, B1 => 
                           REGISTERS_23_63_port, B2 => n407, ZN => n5655);
   U3743 : AOI22_X1 port map( A1 => REGISTERS_17_63_port, A2 => n518, B1 => 
                           REGISTERS_19_63_port, B2 => n481, ZN => n5654);
   U3744 : AOI22_X1 port map( A1 => REGISTERS_20_63_port, A2 => n592, B1 => 
                           REGISTERS_22_63_port, B2 => n555, ZN => n5653);
   U3745 : AOI22_X1 port map( A1 => REGISTERS_16_63_port, A2 => n666, B1 => 
                           REGISTERS_18_63_port, B2 => n629, ZN => n5652);
   U3746 : AND4_X1 port map( A1 => n5655, A2 => n5654, A3 => n5653, A4 => n5652
                           , ZN => n5674);
   U3747 : AOI22_X1 port map( A1 => REGISTERS_29_63_port, A2 => n444, B1 => 
                           REGISTERS_31_63_port, B2 => n407, ZN => n5659);
   U3748 : AOI22_X1 port map( A1 => REGISTERS_25_63_port, A2 => n518, B1 => 
                           REGISTERS_27_63_port, B2 => n481, ZN => n5658);
   U3749 : AOI22_X1 port map( A1 => REGISTERS_28_63_port, A2 => n592, B1 => 
                           REGISTERS_30_63_port, B2 => n555, ZN => n5657);
   U3750 : AOI22_X1 port map( A1 => REGISTERS_24_63_port, A2 => n666, B1 => 
                           REGISTERS_26_63_port, B2 => n629, ZN => n5656);
   U3751 : AND4_X1 port map( A1 => n5659, A2 => n5658, A3 => n5657, A4 => n5656
                           , ZN => n5672);
   U3752 : AOI22_X1 port map( A1 => REGISTERS_5_63_port, A2 => n444, B1 => 
                           REGISTERS_7_63_port, B2 => n407, ZN => n5663);
   U3753 : AOI22_X1 port map( A1 => REGISTERS_1_63_port, A2 => n518, B1 => 
                           REGISTERS_3_63_port, B2 => n481, ZN => n5662);
   U3754 : AOI22_X1 port map( A1 => REGISTERS_4_63_port, A2 => n592, B1 => 
                           REGISTERS_6_63_port, B2 => n555, ZN => n5661);
   U3755 : AOI22_X1 port map( A1 => REGISTERS_0_63_port, A2 => n666, B1 => 
                           REGISTERS_2_63_port, B2 => n629, ZN => n5660);
   U3756 : NAND4_X1 port map( A1 => n5663, A2 => n5662, A3 => n5661, A4 => 
                           n5660, ZN => n5669);
   U3757 : AOI22_X1 port map( A1 => REGISTERS_13_63_port, A2 => n444, B1 => 
                           REGISTERS_15_63_port, B2 => n407, ZN => n5667);
   U3758 : AOI22_X1 port map( A1 => REGISTERS_9_63_port, A2 => n518, B1 => 
                           REGISTERS_11_63_port, B2 => n481, ZN => n5666);
   U3759 : AOI22_X1 port map( A1 => REGISTERS_12_63_port, A2 => n592, B1 => 
                           REGISTERS_14_63_port, B2 => n555, ZN => n5665);
   U3760 : AOI22_X1 port map( A1 => REGISTERS_8_63_port, A2 => n666, B1 => 
                           REGISTERS_10_63_port, B2 => n629, ZN => n5664);
   U3761 : NAND4_X1 port map( A1 => n5667, A2 => n5666, A3 => n5665, A4 => 
                           n5664, ZN => n5668);
   U3762 : AOI22_X1 port map( A1 => n23, A2 => n5669, B1 => n22, B2 => n5668, 
                           ZN => n5670);
   U3763 : OAI221_X1 port map( B1 => n5674, B2 => n5673, C1 => n5672, C2 => 
                           n5671, A => n5670, ZN => N225);
   U3764 : OAI21_X1 port map( B1 => n5924, B2 => n687, A => n5679, ZN => n6052)
                           ;
   U3765 : NAND2_X1 port map( A1 => N288, A2 => n5680, ZN => n5679);
   U3766 : OAI21_X1 port map( B1 => n5925, B2 => n682, A => n5681, ZN => n6053)
                           ;
   U3767 : NAND2_X1 port map( A1 => N287, A2 => n5680, ZN => n5681);
   U3768 : OAI21_X1 port map( B1 => n5926, B2 => n682, A => n5682, ZN => n6054)
                           ;
   U3769 : NAND2_X1 port map( A1 => N286, A2 => n5680, ZN => n5682);
   U3770 : OAI21_X1 port map( B1 => n5927, B2 => n682, A => n5683, ZN => n6055)
                           ;
   U3771 : NAND2_X1 port map( A1 => N285, A2 => n5680, ZN => n5683);
   U3772 : OAI21_X1 port map( B1 => n5928, B2 => n682, A => n5684, ZN => n6056)
                           ;
   U3773 : NAND2_X1 port map( A1 => N284, A2 => n5680, ZN => n5684);
   U3774 : OAI21_X1 port map( B1 => n5929, B2 => n682, A => n5685, ZN => n6057)
                           ;
   U3775 : NAND2_X1 port map( A1 => N283, A2 => n5680, ZN => n5685);
   U3776 : OAI21_X1 port map( B1 => n5930, B2 => n682, A => n5686, ZN => n6058)
                           ;
   U3777 : NAND2_X1 port map( A1 => N282, A2 => n5680, ZN => n5686);
   U3778 : OAI21_X1 port map( B1 => n5931, B2 => n682, A => n5687, ZN => n6059)
                           ;
   U3779 : NAND2_X1 port map( A1 => N281, A2 => n5680, ZN => n5687);
   U3780 : OAI21_X1 port map( B1 => n5932, B2 => n682, A => n5688, ZN => n6060)
                           ;
   U3781 : NAND2_X1 port map( A1 => N280, A2 => n5680, ZN => n5688);
   U3782 : OAI21_X1 port map( B1 => n5933, B2 => n682, A => n5689, ZN => n6061)
                           ;
   U3783 : NAND2_X1 port map( A1 => N279, A2 => n5680, ZN => n5689);
   U3784 : OAI21_X1 port map( B1 => n5934, B2 => n682, A => n5690, ZN => n6062)
                           ;
   U3785 : NAND2_X1 port map( A1 => N278, A2 => n5680, ZN => n5690);
   U3786 : OAI21_X1 port map( B1 => n5935, B2 => n682, A => n5691, ZN => n6063)
                           ;
   U3787 : NAND2_X1 port map( A1 => N277, A2 => n5680, ZN => n5691);
   U3788 : OAI21_X1 port map( B1 => n5936, B2 => n682, A => n5692, ZN => n6064)
                           ;
   U3789 : NAND2_X1 port map( A1 => N276, A2 => n5680, ZN => n5692);
   U3790 : OAI21_X1 port map( B1 => n5937, B2 => n683, A => n5693, ZN => n6065)
                           ;
   U3791 : NAND2_X1 port map( A1 => N275, A2 => n5680, ZN => n5693);
   U3792 : OAI21_X1 port map( B1 => n5938, B2 => n683, A => n5694, ZN => n6066)
                           ;
   U3793 : NAND2_X1 port map( A1 => N274, A2 => n5680, ZN => n5694);
   U3794 : OAI21_X1 port map( B1 => n5939, B2 => n683, A => n5695, ZN => n6067)
                           ;
   U3795 : NAND2_X1 port map( A1 => N273, A2 => n5680, ZN => n5695);
   U3796 : OAI21_X1 port map( B1 => n5940, B2 => n683, A => n5696, ZN => n6068)
                           ;
   U3797 : NAND2_X1 port map( A1 => N272, A2 => n5680, ZN => n5696);
   U3798 : OAI21_X1 port map( B1 => n5941, B2 => n683, A => n5697, ZN => n6069)
                           ;
   U3799 : NAND2_X1 port map( A1 => N271, A2 => n5680, ZN => n5697);
   U3800 : OAI21_X1 port map( B1 => n5942, B2 => n683, A => n5698, ZN => n6070)
                           ;
   U3801 : NAND2_X1 port map( A1 => N270, A2 => n5680, ZN => n5698);
   U3802 : OAI21_X1 port map( B1 => n5943, B2 => n683, A => n5699, ZN => n6071)
                           ;
   U3803 : NAND2_X1 port map( A1 => N269, A2 => n5680, ZN => n5699);
   U3804 : OAI21_X1 port map( B1 => n5944, B2 => n683, A => n5700, ZN => n6072)
                           ;
   U3805 : NAND2_X1 port map( A1 => N268, A2 => n5680, ZN => n5700);
   U3806 : OAI21_X1 port map( B1 => n5945, B2 => n683, A => n5701, ZN => n6073)
                           ;
   U3807 : NAND2_X1 port map( A1 => N267, A2 => n5680, ZN => n5701);
   U3808 : OAI21_X1 port map( B1 => n5946, B2 => n683, A => n5702, ZN => n6074)
                           ;
   U3809 : NAND2_X1 port map( A1 => N266, A2 => n5680, ZN => n5702);
   U3810 : OAI21_X1 port map( B1 => n5947, B2 => n683, A => n5703, ZN => n6075)
                           ;
   U3811 : NAND2_X1 port map( A1 => N265, A2 => n5680, ZN => n5703);
   U3812 : OAI21_X1 port map( B1 => n5948, B2 => n683, A => n5704, ZN => n6076)
                           ;
   U3813 : NAND2_X1 port map( A1 => N264, A2 => n5680, ZN => n5704);
   U3814 : OAI21_X1 port map( B1 => n5949, B2 => n684, A => n5705, ZN => n6077)
                           ;
   U3815 : NAND2_X1 port map( A1 => N263, A2 => n5680, ZN => n5705);
   U3816 : OAI21_X1 port map( B1 => n5950, B2 => n684, A => n5706, ZN => n6078)
                           ;
   U3817 : NAND2_X1 port map( A1 => N262, A2 => n5680, ZN => n5706);
   U3818 : OAI21_X1 port map( B1 => n5951, B2 => n684, A => n5707, ZN => n6079)
                           ;
   U3819 : NAND2_X1 port map( A1 => N261, A2 => n5680, ZN => n5707);
   U3820 : OAI21_X1 port map( B1 => n5952, B2 => n684, A => n5708, ZN => n6080)
                           ;
   U3821 : NAND2_X1 port map( A1 => N260, A2 => n5680, ZN => n5708);
   U3822 : OAI21_X1 port map( B1 => n5953, B2 => n684, A => n5709, ZN => n6081)
                           ;
   U3823 : NAND2_X1 port map( A1 => N259, A2 => n5680, ZN => n5709);
   U3824 : OAI21_X1 port map( B1 => n5954, B2 => n684, A => n5710, ZN => n6082)
                           ;
   U3825 : NAND2_X1 port map( A1 => N258, A2 => n5680, ZN => n5710);
   U3826 : OAI21_X1 port map( B1 => n5955, B2 => n684, A => n5711, ZN => n6083)
                           ;
   U3827 : NAND2_X1 port map( A1 => N257, A2 => n5680, ZN => n5711);
   U3828 : OAI21_X1 port map( B1 => n5956, B2 => n684, A => n5712, ZN => n6084)
                           ;
   U3829 : NAND2_X1 port map( A1 => N256, A2 => n5680, ZN => n5712);
   U3830 : OAI21_X1 port map( B1 => n5957, B2 => n684, A => n5713, ZN => n6085)
                           ;
   U3831 : NAND2_X1 port map( A1 => N255, A2 => n5680, ZN => n5713);
   U3832 : OAI21_X1 port map( B1 => n5958, B2 => n684, A => n5714, ZN => n6086)
                           ;
   U3833 : NAND2_X1 port map( A1 => N254, A2 => n5680, ZN => n5714);
   U3834 : OAI21_X1 port map( B1 => n5959, B2 => n684, A => n5715, ZN => n6087)
                           ;
   U3835 : NAND2_X1 port map( A1 => N253, A2 => n5680, ZN => n5715);
   U3836 : OAI21_X1 port map( B1 => n5960, B2 => n684, A => n5716, ZN => n6088)
                           ;
   U3837 : NAND2_X1 port map( A1 => N252, A2 => n5680, ZN => n5716);
   U3838 : OAI21_X1 port map( B1 => n5961, B2 => n685, A => n5717, ZN => n6089)
                           ;
   U3839 : NAND2_X1 port map( A1 => N251, A2 => n5680, ZN => n5717);
   U3840 : OAI21_X1 port map( B1 => n5962, B2 => n685, A => n5718, ZN => n6090)
                           ;
   U3841 : NAND2_X1 port map( A1 => N250, A2 => n5680, ZN => n5718);
   U3842 : OAI21_X1 port map( B1 => n5963, B2 => n685, A => n5719, ZN => n6091)
                           ;
   U3843 : NAND2_X1 port map( A1 => N249, A2 => n5680, ZN => n5719);
   U3844 : OAI21_X1 port map( B1 => n5964, B2 => n685, A => n5720, ZN => n6092)
                           ;
   U3845 : NAND2_X1 port map( A1 => N248, A2 => n5680, ZN => n5720);
   U3846 : OAI21_X1 port map( B1 => n5965, B2 => n685, A => n5721, ZN => n6093)
                           ;
   U3847 : NAND2_X1 port map( A1 => N247, A2 => n5680, ZN => n5721);
   U3848 : OAI21_X1 port map( B1 => n5966, B2 => n685, A => n5722, ZN => n6094)
                           ;
   U3849 : NAND2_X1 port map( A1 => N246, A2 => n5680, ZN => n5722);
   U3850 : OAI21_X1 port map( B1 => n5967, B2 => n685, A => n5723, ZN => n6095)
                           ;
   U3851 : NAND2_X1 port map( A1 => N245, A2 => n5680, ZN => n5723);
   U3852 : OAI21_X1 port map( B1 => n5968, B2 => n685, A => n5724, ZN => n6096)
                           ;
   U3853 : NAND2_X1 port map( A1 => N244, A2 => n5680, ZN => n5724);
   U3854 : OAI21_X1 port map( B1 => n5969, B2 => n685, A => n5725, ZN => n6097)
                           ;
   U3855 : NAND2_X1 port map( A1 => N243, A2 => n5680, ZN => n5725);
   U3856 : OAI21_X1 port map( B1 => n5970, B2 => n685, A => n5726, ZN => n6098)
                           ;
   U3857 : NAND2_X1 port map( A1 => N242, A2 => n5680, ZN => n5726);
   U3858 : OAI21_X1 port map( B1 => n5971, B2 => n685, A => n5727, ZN => n6099)
                           ;
   U3859 : NAND2_X1 port map( A1 => N241, A2 => n5680, ZN => n5727);
   U3860 : OAI21_X1 port map( B1 => n5972, B2 => n685, A => n5728, ZN => n6100)
                           ;
   U3861 : NAND2_X1 port map( A1 => N240, A2 => n5680, ZN => n5728);
   U3862 : OAI21_X1 port map( B1 => n5973, B2 => n686, A => n5729, ZN => n6101)
                           ;
   U3863 : NAND2_X1 port map( A1 => N239, A2 => n5680, ZN => n5729);
   U3864 : OAI21_X1 port map( B1 => n5974, B2 => n686, A => n5730, ZN => n6102)
                           ;
   U3865 : NAND2_X1 port map( A1 => N238, A2 => n5680, ZN => n5730);
   U3866 : OAI21_X1 port map( B1 => n5975, B2 => n686, A => n5731, ZN => n6103)
                           ;
   U3867 : NAND2_X1 port map( A1 => N237, A2 => n5680, ZN => n5731);
   U3868 : OAI21_X1 port map( B1 => n5976, B2 => n686, A => n5732, ZN => n6104)
                           ;
   U3869 : NAND2_X1 port map( A1 => N236, A2 => n5680, ZN => n5732);
   U3870 : OAI21_X1 port map( B1 => n5977, B2 => n686, A => n5733, ZN => n6105)
                           ;
   U3871 : NAND2_X1 port map( A1 => N235, A2 => n5680, ZN => n5733);
   U3872 : OAI21_X1 port map( B1 => n5978, B2 => n686, A => n5734, ZN => n6106)
                           ;
   U3873 : NAND2_X1 port map( A1 => N234, A2 => n5680, ZN => n5734);
   U3874 : OAI21_X1 port map( B1 => n5979, B2 => n686, A => n5735, ZN => n6107)
                           ;
   U3875 : NAND2_X1 port map( A1 => N233, A2 => n5680, ZN => n5735);
   U3876 : OAI21_X1 port map( B1 => n5980, B2 => n686, A => n5736, ZN => n6108)
                           ;
   U3877 : NAND2_X1 port map( A1 => N232, A2 => n5680, ZN => n5736);
   U3878 : OAI21_X1 port map( B1 => n5981, B2 => n686, A => n5737, ZN => n6109)
                           ;
   U3879 : NAND2_X1 port map( A1 => N231, A2 => n5680, ZN => n5737);
   U3880 : OAI21_X1 port map( B1 => n5982, B2 => n686, A => n5738, ZN => n6110)
                           ;
   U3881 : NAND2_X1 port map( A1 => N230, A2 => n5680, ZN => n5738);
   U3882 : OAI21_X1 port map( B1 => n5983, B2 => n686, A => n5739, ZN => n6111)
                           ;
   U3883 : NAND2_X1 port map( A1 => N229, A2 => n5680, ZN => n5739);
   U3884 : OAI21_X1 port map( B1 => n5984, B2 => n686, A => n5740, ZN => n6112)
                           ;
   U3885 : NAND2_X1 port map( A1 => N228, A2 => n5680, ZN => n5740);
   U3886 : OAI21_X1 port map( B1 => n5985, B2 => n687, A => n5741, ZN => n6113)
                           ;
   U3887 : NAND2_X1 port map( A1 => N227, A2 => n5680, ZN => n5741);
   U3888 : OAI21_X1 port map( B1 => n5986, B2 => n687, A => n5742, ZN => n6114)
                           ;
   U3889 : NAND2_X1 port map( A1 => N226, A2 => n5680, ZN => n5742);
   U3890 : OAI21_X1 port map( B1 => n5987, B2 => n687, A => n5743, ZN => n6115)
                           ;
   U3891 : NAND2_X1 port map( A1 => N225, A2 => n5680, ZN => n5743);
   U3892 : OAI21_X1 port map( B1 => n5988, B2 => n687, A => n5745, ZN => n6116)
                           ;
   U3893 : NAND2_X1 port map( A1 => N159, A2 => n5746, ZN => n5745);
   U3894 : OAI21_X1 port map( B1 => n5989, B2 => n687, A => n5747, ZN => n6117)
                           ;
   U3895 : NAND2_X1 port map( A1 => N158, A2 => n5746, ZN => n5747);
   U3896 : OAI21_X1 port map( B1 => n5990, B2 => n687, A => n5748, ZN => n6118)
                           ;
   U3897 : NAND2_X1 port map( A1 => N157, A2 => n5746, ZN => n5748);
   U3898 : OAI21_X1 port map( B1 => n5991, B2 => n687, A => n5749, ZN => n6119)
                           ;
   U3899 : NAND2_X1 port map( A1 => N156, A2 => n5746, ZN => n5749);
   U3900 : OAI21_X1 port map( B1 => n5992, B2 => n687, A => n5750, ZN => n6120)
                           ;
   U3901 : NAND2_X1 port map( A1 => N155, A2 => n5746, ZN => n5750);
   U3902 : OAI21_X1 port map( B1 => n5993, B2 => n687, A => n5751, ZN => n6121)
                           ;
   U3903 : NAND2_X1 port map( A1 => N154, A2 => n5746, ZN => n5751);
   U3904 : OAI21_X1 port map( B1 => n5994, B2 => n687, A => n5752, ZN => n6122)
                           ;
   U3905 : NAND2_X1 port map( A1 => N153, A2 => n5746, ZN => n5752);
   U3906 : OAI21_X1 port map( B1 => n5995, B2 => n688, A => n5753, ZN => n6123)
                           ;
   U3907 : NAND2_X1 port map( A1 => N152, A2 => n5746, ZN => n5753);
   U3908 : OAI21_X1 port map( B1 => n5996, B2 => n687, A => n5754, ZN => n6124)
                           ;
   U3909 : NAND2_X1 port map( A1 => N151, A2 => n5746, ZN => n5754);
   U3910 : OAI21_X1 port map( B1 => n5997, B2 => n688, A => n5755, ZN => n6125)
                           ;
   U3911 : NAND2_X1 port map( A1 => N150, A2 => n5746, ZN => n5755);
   U3912 : OAI21_X1 port map( B1 => n5998, B2 => n688, A => n5756, ZN => n6126)
                           ;
   U3913 : NAND2_X1 port map( A1 => N149, A2 => n5746, ZN => n5756);
   U3914 : OAI21_X1 port map( B1 => n5999, B2 => n688, A => n5757, ZN => n6127)
                           ;
   U3915 : NAND2_X1 port map( A1 => N148, A2 => n5746, ZN => n5757);
   U3916 : OAI21_X1 port map( B1 => n6000, B2 => n688, A => n5758, ZN => n6128)
                           ;
   U3917 : NAND2_X1 port map( A1 => N147, A2 => n5746, ZN => n5758);
   U3918 : OAI21_X1 port map( B1 => n6001, B2 => n688, A => n5759, ZN => n6129)
                           ;
   U3919 : NAND2_X1 port map( A1 => N146, A2 => n5746, ZN => n5759);
   U3920 : OAI21_X1 port map( B1 => n6002, B2 => n688, A => n5760, ZN => n6130)
                           ;
   U3921 : NAND2_X1 port map( A1 => N145, A2 => n5746, ZN => n5760);
   U3922 : OAI21_X1 port map( B1 => n6003, B2 => n688, A => n5761, ZN => n6131)
                           ;
   U3923 : NAND2_X1 port map( A1 => N144, A2 => n5746, ZN => n5761);
   U3924 : OAI21_X1 port map( B1 => n6004, B2 => n688, A => n5762, ZN => n6132)
                           ;
   U3925 : NAND2_X1 port map( A1 => N143, A2 => n5746, ZN => n5762);
   U3926 : OAI21_X1 port map( B1 => n6005, B2 => n688, A => n5763, ZN => n6133)
                           ;
   U3927 : NAND2_X1 port map( A1 => N142, A2 => n5746, ZN => n5763);
   U3928 : OAI21_X1 port map( B1 => n6006, B2 => n688, A => n5764, ZN => n6134)
                           ;
   U3929 : NAND2_X1 port map( A1 => N141, A2 => n5746, ZN => n5764);
   U3930 : OAI21_X1 port map( B1 => n6007, B2 => n689, A => n5765, ZN => n6135)
                           ;
   U3931 : NAND2_X1 port map( A1 => N140, A2 => n5746, ZN => n5765);
   U3932 : OAI21_X1 port map( B1 => n6008, B2 => n688, A => n5766, ZN => n6136)
                           ;
   U3933 : NAND2_X1 port map( A1 => N139, A2 => n5746, ZN => n5766);
   U3934 : OAI21_X1 port map( B1 => n6009, B2 => n689, A => n5767, ZN => n6137)
                           ;
   U3935 : NAND2_X1 port map( A1 => N138, A2 => n5746, ZN => n5767);
   U3936 : OAI21_X1 port map( B1 => n6010, B2 => n689, A => n5768, ZN => n6138)
                           ;
   U3937 : NAND2_X1 port map( A1 => N137, A2 => n5746, ZN => n5768);
   U3938 : OAI21_X1 port map( B1 => n6011, B2 => n689, A => n5769, ZN => n6139)
                           ;
   U3939 : NAND2_X1 port map( A1 => N136, A2 => n5746, ZN => n5769);
   U3940 : OAI21_X1 port map( B1 => n6012, B2 => n689, A => n5770, ZN => n6140)
                           ;
   U3941 : NAND2_X1 port map( A1 => N135, A2 => n5746, ZN => n5770);
   U3942 : OAI21_X1 port map( B1 => n6013, B2 => n689, A => n5771, ZN => n6141)
                           ;
   U3943 : NAND2_X1 port map( A1 => N134, A2 => n5746, ZN => n5771);
   U3944 : OAI21_X1 port map( B1 => n6014, B2 => n689, A => n5772, ZN => n6142)
                           ;
   U3945 : NAND2_X1 port map( A1 => N133, A2 => n5746, ZN => n5772);
   U3946 : OAI21_X1 port map( B1 => n6015, B2 => n689, A => n5773, ZN => n6143)
                           ;
   U3947 : NAND2_X1 port map( A1 => N132, A2 => n5746, ZN => n5773);
   U3948 : OAI21_X1 port map( B1 => n6016, B2 => n689, A => n5774, ZN => n6144)
                           ;
   U3949 : NAND2_X1 port map( A1 => N131, A2 => n5746, ZN => n5774);
   U3950 : OAI21_X1 port map( B1 => n6017, B2 => n689, A => n5775, ZN => n6145)
                           ;
   U3951 : NAND2_X1 port map( A1 => N130, A2 => n5746, ZN => n5775);
   U3952 : OAI21_X1 port map( B1 => n6018, B2 => n689, A => n5776, ZN => n6146)
                           ;
   U3953 : NAND2_X1 port map( A1 => N129, A2 => n5746, ZN => n5776);
   U3954 : OAI21_X1 port map( B1 => n6019, B2 => n690, A => n5777, ZN => n6147)
                           ;
   U3955 : NAND2_X1 port map( A1 => N128, A2 => n5746, ZN => n5777);
   U3956 : OAI21_X1 port map( B1 => n6020, B2 => n689, A => n5778, ZN => n6148)
                           ;
   U3957 : NAND2_X1 port map( A1 => N127, A2 => n5746, ZN => n5778);
   U3958 : OAI21_X1 port map( B1 => n6021, B2 => n690, A => n5779, ZN => n6149)
                           ;
   U3959 : NAND2_X1 port map( A1 => N126, A2 => n5746, ZN => n5779);
   U3960 : OAI21_X1 port map( B1 => n6022, B2 => n690, A => n5780, ZN => n6150)
                           ;
   U3961 : NAND2_X1 port map( A1 => N125, A2 => n5746, ZN => n5780);
   U3962 : OAI21_X1 port map( B1 => n6023, B2 => n690, A => n5781, ZN => n6151)
                           ;
   U3963 : NAND2_X1 port map( A1 => N124, A2 => n5746, ZN => n5781);
   U3964 : OAI21_X1 port map( B1 => n6024, B2 => n690, A => n5782, ZN => n6152)
                           ;
   U3965 : NAND2_X1 port map( A1 => N123, A2 => n5746, ZN => n5782);
   U3966 : OAI21_X1 port map( B1 => n6025, B2 => n690, A => n5783, ZN => n6153)
                           ;
   U3967 : NAND2_X1 port map( A1 => N122, A2 => n5746, ZN => n5783);
   U3968 : OAI21_X1 port map( B1 => n6026, B2 => n690, A => n5784, ZN => n6154)
                           ;
   U3969 : NAND2_X1 port map( A1 => N121, A2 => n5746, ZN => n5784);
   U3970 : OAI21_X1 port map( B1 => n6027, B2 => n690, A => n5785, ZN => n6155)
                           ;
   U3971 : NAND2_X1 port map( A1 => N120, A2 => n5746, ZN => n5785);
   U3972 : OAI21_X1 port map( B1 => n6028, B2 => n690, A => n5786, ZN => n6156)
                           ;
   U3973 : NAND2_X1 port map( A1 => N119, A2 => n5746, ZN => n5786);
   U3974 : OAI21_X1 port map( B1 => n6029, B2 => n690, A => n5787, ZN => n6157)
                           ;
   U3975 : NAND2_X1 port map( A1 => N118, A2 => n5746, ZN => n5787);
   U3976 : OAI21_X1 port map( B1 => n6030, B2 => n690, A => n5788, ZN => n6158)
                           ;
   U3977 : NAND2_X1 port map( A1 => N117, A2 => n5746, ZN => n5788);
   U3978 : OAI21_X1 port map( B1 => n6031, B2 => n691, A => n5789, ZN => n6159)
                           ;
   U3979 : NAND2_X1 port map( A1 => N116, A2 => n5746, ZN => n5789);
   U3980 : OAI21_X1 port map( B1 => n6032, B2 => n690, A => n5790, ZN => n6160)
                           ;
   U3981 : NAND2_X1 port map( A1 => N115, A2 => n5746, ZN => n5790);
   U3982 : OAI21_X1 port map( B1 => n6033, B2 => n691, A => n5791, ZN => n6161)
                           ;
   U3983 : NAND2_X1 port map( A1 => N114, A2 => n5746, ZN => n5791);
   U3984 : OAI21_X1 port map( B1 => n6034, B2 => n691, A => n5792, ZN => n6162)
                           ;
   U3985 : NAND2_X1 port map( A1 => N113, A2 => n5746, ZN => n5792);
   U3986 : OAI21_X1 port map( B1 => n6035, B2 => n691, A => n5793, ZN => n6163)
                           ;
   U3987 : NAND2_X1 port map( A1 => N112, A2 => n5746, ZN => n5793);
   U3988 : OAI21_X1 port map( B1 => n6036, B2 => n691, A => n5794, ZN => n6164)
                           ;
   U3989 : NAND2_X1 port map( A1 => N111, A2 => n5746, ZN => n5794);
   U3990 : OAI21_X1 port map( B1 => n6037, B2 => n691, A => n5795, ZN => n6165)
                           ;
   U3991 : NAND2_X1 port map( A1 => N110, A2 => n5746, ZN => n5795);
   U3992 : OAI21_X1 port map( B1 => n6038, B2 => n691, A => n5796, ZN => n6166)
                           ;
   U3993 : NAND2_X1 port map( A1 => N109, A2 => n5746, ZN => n5796);
   U3994 : OAI21_X1 port map( B1 => n6039, B2 => n691, A => n5797, ZN => n6167)
                           ;
   U3995 : NAND2_X1 port map( A1 => N108, A2 => n5746, ZN => n5797);
   U3996 : OAI21_X1 port map( B1 => n6040, B2 => n691, A => n5798, ZN => n6168)
                           ;
   U3997 : NAND2_X1 port map( A1 => N107, A2 => n5746, ZN => n5798);
   U3998 : OAI21_X1 port map( B1 => n6041, B2 => n691, A => n5799, ZN => n6169)
                           ;
   U3999 : NAND2_X1 port map( A1 => N106, A2 => n5746, ZN => n5799);
   U4000 : OAI21_X1 port map( B1 => n6042, B2 => n691, A => n5800, ZN => n6170)
                           ;
   U4001 : NAND2_X1 port map( A1 => N105, A2 => n5746, ZN => n5800);
   U4002 : OAI21_X1 port map( B1 => n6043, B2 => n692, A => n5801, ZN => n6171)
                           ;
   U4003 : NAND2_X1 port map( A1 => N104, A2 => n5746, ZN => n5801);
   U4004 : OAI21_X1 port map( B1 => n6044, B2 => n691, A => n5802, ZN => n6172)
                           ;
   U4005 : NAND2_X1 port map( A1 => N103, A2 => n5746, ZN => n5802);
   U4006 : OAI21_X1 port map( B1 => n6045, B2 => n692, A => n5803, ZN => n6173)
                           ;
   U4007 : NAND2_X1 port map( A1 => N102, A2 => n5746, ZN => n5803);
   U4008 : OAI21_X1 port map( B1 => n6046, B2 => n692, A => n5804, ZN => n6174)
                           ;
   U4009 : NAND2_X1 port map( A1 => N101, A2 => n5746, ZN => n5804);
   U4010 : OAI21_X1 port map( B1 => n6047, B2 => n692, A => n5805, ZN => n6175)
                           ;
   U4011 : NAND2_X1 port map( A1 => N100, A2 => n5746, ZN => n5805);
   U4012 : OAI21_X1 port map( B1 => n6048, B2 => n692, A => n5806, ZN => n6176)
                           ;
   U4013 : NAND2_X1 port map( A1 => N99, A2 => n5746, ZN => n5806);
   U4014 : OAI21_X1 port map( B1 => n6049, B2 => n692, A => n5807, ZN => n6177)
                           ;
   U4015 : NAND2_X1 port map( A1 => N98, A2 => n5746, ZN => n5807);
   U4016 : OAI21_X1 port map( B1 => n6050, B2 => n692, A => n5808, ZN => n6178)
                           ;
   U4017 : NAND2_X1 port map( A1 => N97, A2 => n5746, ZN => n5808);
   U4018 : OAI21_X1 port map( B1 => n6051, B2 => n692, A => n5809, ZN => n6179)
                           ;
   U4019 : NAND2_X1 port map( A1 => N96, A2 => n5746, ZN => n5809);
   U4020 : MUX2_X1 port map( A => REGISTERS_0_63_port, B => n5810, S => n85, Z 
                           => n4503);
   U4021 : MUX2_X1 port map( A => REGISTERS_0_62_port, B => n5812, S => n85, Z 
                           => n4502);
   U4022 : MUX2_X1 port map( A => REGISTERS_0_61_port, B => n5813, S => n85, Z 
                           => n4501);
   U4023 : MUX2_X1 port map( A => REGISTERS_0_60_port, B => n5814, S => n85, Z 
                           => n4500);
   U4024 : MUX2_X1 port map( A => REGISTERS_0_59_port, B => n5815, S => n85, Z 
                           => n4499);
   U4025 : MUX2_X1 port map( A => REGISTERS_0_58_port, B => n5816, S => n85, Z 
                           => n4498);
   U4026 : MUX2_X1 port map( A => REGISTERS_0_57_port, B => n5817, S => n85, Z 
                           => n4497);
   U4027 : MUX2_X1 port map( A => REGISTERS_0_56_port, B => n5818, S => n85, Z 
                           => n4496);
   U4028 : MUX2_X1 port map( A => REGISTERS_0_55_port, B => n5819, S => n85, Z 
                           => n4495);
   U4029 : MUX2_X1 port map( A => REGISTERS_0_54_port, B => n5820, S => n85, Z 
                           => n4494);
   U4030 : MUX2_X1 port map( A => REGISTERS_0_53_port, B => n5821, S => n85, Z 
                           => n4493);
   U4031 : MUX2_X1 port map( A => REGISTERS_0_52_port, B => n5822, S => n85, Z 
                           => n4492);
   U4032 : MUX2_X1 port map( A => REGISTERS_0_51_port, B => n5823, S => n85, Z 
                           => n4491);
   U4033 : MUX2_X1 port map( A => REGISTERS_0_50_port, B => n5824, S => n85, Z 
                           => n4490);
   U4034 : MUX2_X1 port map( A => REGISTERS_0_49_port, B => n5825, S => n85, Z 
                           => n4489);
   U4035 : MUX2_X1 port map( A => REGISTERS_0_48_port, B => n5826, S => n85, Z 
                           => n4488);
   U4036 : MUX2_X1 port map( A => REGISTERS_0_47_port, B => n5827, S => n85, Z 
                           => n4487);
   U4037 : MUX2_X1 port map( A => REGISTERS_0_46_port, B => n5828, S => n85, Z 
                           => n4486);
   U4038 : MUX2_X1 port map( A => REGISTERS_0_45_port, B => n5829, S => n85, Z 
                           => n4485);
   U4039 : MUX2_X1 port map( A => REGISTERS_0_44_port, B => n5830, S => n85, Z 
                           => n4484);
   U4040 : MUX2_X1 port map( A => REGISTERS_0_43_port, B => n5831, S => n85, Z 
                           => n4483);
   U4041 : MUX2_X1 port map( A => REGISTERS_0_42_port, B => n5832, S => n85, Z 
                           => n4482);
   U4042 : MUX2_X1 port map( A => REGISTERS_0_41_port, B => n5833, S => n85, Z 
                           => n4481);
   U4043 : MUX2_X1 port map( A => REGISTERS_0_40_port, B => n5834, S => n85, Z 
                           => n4480);
   U4044 : MUX2_X1 port map( A => REGISTERS_0_39_port, B => n5835, S => n85, Z 
                           => n4479);
   U4045 : MUX2_X1 port map( A => REGISTERS_0_38_port, B => n5836, S => n85, Z 
                           => n4478);
   U4046 : MUX2_X1 port map( A => REGISTERS_0_37_port, B => n5837, S => n85, Z 
                           => n4477);
   U4047 : MUX2_X1 port map( A => REGISTERS_0_36_port, B => n5838, S => n85, Z 
                           => n4476);
   U4048 : MUX2_X1 port map( A => REGISTERS_0_35_port, B => n5839, S => n85, Z 
                           => n4475);
   U4049 : MUX2_X1 port map( A => REGISTERS_0_34_port, B => n5840, S => n85, Z 
                           => n4474);
   U4050 : MUX2_X1 port map( A => REGISTERS_0_33_port, B => n5841, S => n85, Z 
                           => n4473);
   U4051 : MUX2_X1 port map( A => REGISTERS_0_32_port, B => n5842, S => n85, Z 
                           => n4472);
   U4052 : MUX2_X1 port map( A => REGISTERS_0_31_port, B => n5843, S => n85, Z 
                           => n4471);
   U4053 : MUX2_X1 port map( A => REGISTERS_0_30_port, B => n5844, S => n85, Z 
                           => n4470);
   U4054 : MUX2_X1 port map( A => REGISTERS_0_29_port, B => n5845, S => n85, Z 
                           => n4469);
   U4055 : MUX2_X1 port map( A => REGISTERS_0_28_port, B => n5846, S => n85, Z 
                           => n4468);
   U4056 : MUX2_X1 port map( A => REGISTERS_0_27_port, B => n5847, S => n85, Z 
                           => n4467);
   U4057 : MUX2_X1 port map( A => REGISTERS_0_26_port, B => n5848, S => n85, Z 
                           => n4466);
   U4058 : MUX2_X1 port map( A => REGISTERS_0_25_port, B => n5849, S => n85, Z 
                           => n4465);
   U4059 : MUX2_X1 port map( A => REGISTERS_0_24_port, B => n5850, S => n85, Z 
                           => n4464);
   U4060 : MUX2_X1 port map( A => REGISTERS_0_23_port, B => n5851, S => n85, Z 
                           => n4463);
   U4061 : MUX2_X1 port map( A => REGISTERS_0_22_port, B => n5852, S => n85, Z 
                           => n4462);
   U4062 : MUX2_X1 port map( A => REGISTERS_0_21_port, B => n5853, S => n85, Z 
                           => n4461);
   U4063 : MUX2_X1 port map( A => REGISTERS_0_20_port, B => n5854, S => n85, Z 
                           => n4460);
   U4064 : MUX2_X1 port map( A => REGISTERS_0_19_port, B => n5855, S => n85, Z 
                           => n4459);
   U4065 : MUX2_X1 port map( A => REGISTERS_0_18_port, B => n5856, S => n85, Z 
                           => n4458);
   U4066 : MUX2_X1 port map( A => REGISTERS_0_17_port, B => n5857, S => n85, Z 
                           => n4457);
   U4067 : MUX2_X1 port map( A => REGISTERS_0_16_port, B => n5858, S => n85, Z 
                           => n4456);
   U4068 : MUX2_X1 port map( A => REGISTERS_0_15_port, B => n5859, S => n85, Z 
                           => n4455);
   U4069 : MUX2_X1 port map( A => REGISTERS_0_14_port, B => n5860, S => n85, Z 
                           => n4454);
   U4070 : MUX2_X1 port map( A => REGISTERS_0_13_port, B => n5861, S => n85, Z 
                           => n4453);
   U4071 : MUX2_X1 port map( A => REGISTERS_0_12_port, B => n5862, S => n85, Z 
                           => n4452);
   U4072 : MUX2_X1 port map( A => REGISTERS_0_11_port, B => n5863, S => n85, Z 
                           => n4451);
   U4073 : MUX2_X1 port map( A => REGISTERS_0_10_port, B => n5864, S => n85, Z 
                           => n4450);
   U4074 : MUX2_X1 port map( A => REGISTERS_0_9_port, B => n5865, S => n85, Z 
                           => n4449);
   U4075 : MUX2_X1 port map( A => REGISTERS_0_8_port, B => n5866, S => n85, Z 
                           => n4448);
   U4076 : MUX2_X1 port map( A => REGISTERS_0_7_port, B => n5867, S => n85, Z 
                           => n4447);
   U4077 : MUX2_X1 port map( A => REGISTERS_0_6_port, B => n5868, S => n85, Z 
                           => n4446);
   U4078 : MUX2_X1 port map( A => REGISTERS_0_5_port, B => n5869, S => n85, Z 
                           => n4445);
   U4079 : MUX2_X1 port map( A => REGISTERS_0_4_port, B => n5870, S => n85, Z 
                           => n4444);
   U4080 : MUX2_X1 port map( A => REGISTERS_0_3_port, B => n5871, S => n85, Z 
                           => n4443);
   U4081 : MUX2_X1 port map( A => REGISTERS_0_2_port, B => n5872, S => n85, Z 
                           => n4442);
   U4082 : MUX2_X1 port map( A => REGISTERS_0_1_port, B => n5873, S => n85, Z 
                           => n4441);
   U4083 : MUX2_X1 port map( A => REGISTERS_0_0_port, B => n5874, S => n85, Z 
                           => n4440);
   U4084 : OAI21_X1 port map( B1 => n5875, B2 => n5876, A => n5744, ZN => n5811
                           );
   U4085 : MUX2_X1 port map( A => REGISTERS_1_63_port, B => n5810, S => n87, Z 
                           => n4439);
   U4086 : MUX2_X1 port map( A => REGISTERS_1_62_port, B => n5812, S => n87, Z 
                           => n4438);
   U4087 : MUX2_X1 port map( A => REGISTERS_1_61_port, B => n5813, S => n87, Z 
                           => n4437);
   U4088 : MUX2_X1 port map( A => REGISTERS_1_60_port, B => n5814, S => n87, Z 
                           => n4436);
   U4089 : MUX2_X1 port map( A => REGISTERS_1_59_port, B => n5815, S => n87, Z 
                           => n4435);
   U4090 : MUX2_X1 port map( A => REGISTERS_1_58_port, B => n5816, S => n87, Z 
                           => n4434);
   U4091 : MUX2_X1 port map( A => REGISTERS_1_57_port, B => n5817, S => n87, Z 
                           => n4433);
   U4092 : MUX2_X1 port map( A => REGISTERS_1_56_port, B => n5818, S => n87, Z 
                           => n4432);
   U4093 : MUX2_X1 port map( A => REGISTERS_1_55_port, B => n5819, S => n87, Z 
                           => n4431);
   U4094 : MUX2_X1 port map( A => REGISTERS_1_54_port, B => n5820, S => n87, Z 
                           => n4430);
   U4095 : MUX2_X1 port map( A => REGISTERS_1_53_port, B => n5821, S => n87, Z 
                           => n4429);
   U4096 : MUX2_X1 port map( A => REGISTERS_1_52_port, B => n5822, S => n87, Z 
                           => n4428);
   U4097 : MUX2_X1 port map( A => REGISTERS_1_51_port, B => n5823, S => n87, Z 
                           => n4427);
   U4098 : MUX2_X1 port map( A => REGISTERS_1_50_port, B => n5824, S => n87, Z 
                           => n4426);
   U4099 : MUX2_X1 port map( A => REGISTERS_1_49_port, B => n5825, S => n87, Z 
                           => n4425);
   U4100 : MUX2_X1 port map( A => REGISTERS_1_48_port, B => n5826, S => n87, Z 
                           => n4424);
   U4101 : MUX2_X1 port map( A => REGISTERS_1_47_port, B => n5827, S => n87, Z 
                           => n4423);
   U4102 : MUX2_X1 port map( A => REGISTERS_1_46_port, B => n5828, S => n87, Z 
                           => n4422);
   U4103 : MUX2_X1 port map( A => REGISTERS_1_45_port, B => n5829, S => n87, Z 
                           => n4421);
   U4104 : MUX2_X1 port map( A => REGISTERS_1_44_port, B => n5830, S => n87, Z 
                           => n4420);
   U4105 : MUX2_X1 port map( A => REGISTERS_1_43_port, B => n5831, S => n87, Z 
                           => n4419);
   U4106 : MUX2_X1 port map( A => REGISTERS_1_42_port, B => n5832, S => n87, Z 
                           => n4418);
   U4107 : MUX2_X1 port map( A => REGISTERS_1_41_port, B => n5833, S => n87, Z 
                           => n4417);
   U4108 : MUX2_X1 port map( A => REGISTERS_1_40_port, B => n5834, S => n87, Z 
                           => n4416);
   U4109 : MUX2_X1 port map( A => REGISTERS_1_39_port, B => n5835, S => n87, Z 
                           => n4415);
   U4110 : MUX2_X1 port map( A => REGISTERS_1_38_port, B => n5836, S => n87, Z 
                           => n4414);
   U4111 : MUX2_X1 port map( A => REGISTERS_1_37_port, B => n5837, S => n87, Z 
                           => n4413);
   U4112 : MUX2_X1 port map( A => REGISTERS_1_36_port, B => n5838, S => n87, Z 
                           => n4412);
   U4113 : MUX2_X1 port map( A => REGISTERS_1_35_port, B => n5839, S => n87, Z 
                           => n4411);
   U4114 : MUX2_X1 port map( A => REGISTERS_1_34_port, B => n5840, S => n87, Z 
                           => n4410);
   U4115 : MUX2_X1 port map( A => REGISTERS_1_33_port, B => n5841, S => n87, Z 
                           => n4409);
   U4116 : MUX2_X1 port map( A => REGISTERS_1_32_port, B => n5842, S => n87, Z 
                           => n4408);
   U4117 : MUX2_X1 port map( A => REGISTERS_1_31_port, B => n5843, S => n87, Z 
                           => n4407);
   U4118 : MUX2_X1 port map( A => REGISTERS_1_30_port, B => n5844, S => n87, Z 
                           => n4406);
   U4119 : MUX2_X1 port map( A => REGISTERS_1_29_port, B => n5845, S => n87, Z 
                           => n4405);
   U4120 : MUX2_X1 port map( A => REGISTERS_1_28_port, B => n5846, S => n87, Z 
                           => n4404);
   U4121 : MUX2_X1 port map( A => REGISTERS_1_27_port, B => n5847, S => n87, Z 
                           => n4403);
   U4122 : MUX2_X1 port map( A => REGISTERS_1_26_port, B => n5848, S => n87, Z 
                           => n4402);
   U4123 : MUX2_X1 port map( A => REGISTERS_1_25_port, B => n5849, S => n87, Z 
                           => n4401);
   U4124 : MUX2_X1 port map( A => REGISTERS_1_24_port, B => n5850, S => n87, Z 
                           => n4400);
   U4125 : MUX2_X1 port map( A => REGISTERS_1_23_port, B => n5851, S => n87, Z 
                           => n4399);
   U4126 : MUX2_X1 port map( A => REGISTERS_1_22_port, B => n5852, S => n87, Z 
                           => n4398);
   U4127 : MUX2_X1 port map( A => REGISTERS_1_21_port, B => n5853, S => n87, Z 
                           => n4397);
   U4128 : MUX2_X1 port map( A => REGISTERS_1_20_port, B => n5854, S => n87, Z 
                           => n4396);
   U4129 : MUX2_X1 port map( A => REGISTERS_1_19_port, B => n5855, S => n87, Z 
                           => n4395);
   U4130 : MUX2_X1 port map( A => REGISTERS_1_18_port, B => n5856, S => n87, Z 
                           => n4394);
   U4131 : MUX2_X1 port map( A => REGISTERS_1_17_port, B => n5857, S => n87, Z 
                           => n4393);
   U4132 : MUX2_X1 port map( A => REGISTERS_1_16_port, B => n5858, S => n87, Z 
                           => n4392);
   U4133 : MUX2_X1 port map( A => REGISTERS_1_15_port, B => n5859, S => n87, Z 
                           => n4391);
   U4134 : MUX2_X1 port map( A => REGISTERS_1_14_port, B => n5860, S => n87, Z 
                           => n4390);
   U4135 : MUX2_X1 port map( A => REGISTERS_1_13_port, B => n5861, S => n87, Z 
                           => n4389);
   U4136 : MUX2_X1 port map( A => REGISTERS_1_12_port, B => n5862, S => n87, Z 
                           => n4388);
   U4137 : MUX2_X1 port map( A => REGISTERS_1_11_port, B => n5863, S => n87, Z 
                           => n4387);
   U4138 : MUX2_X1 port map( A => REGISTERS_1_10_port, B => n5864, S => n87, Z 
                           => n4386);
   U4139 : MUX2_X1 port map( A => REGISTERS_1_9_port, B => n5865, S => n87, Z 
                           => n4385);
   U4140 : MUX2_X1 port map( A => REGISTERS_1_8_port, B => n5866, S => n87, Z 
                           => n4384);
   U4141 : MUX2_X1 port map( A => REGISTERS_1_7_port, B => n5867, S => n87, Z 
                           => n4383);
   U4142 : MUX2_X1 port map( A => REGISTERS_1_6_port, B => n5868, S => n87, Z 
                           => n4382);
   U4143 : MUX2_X1 port map( A => REGISTERS_1_5_port, B => n5869, S => n87, Z 
                           => n4381);
   U4144 : MUX2_X1 port map( A => REGISTERS_1_4_port, B => n5870, S => n87, Z 
                           => n4380);
   U4145 : MUX2_X1 port map( A => REGISTERS_1_3_port, B => n5871, S => n87, Z 
                           => n4379);
   U4146 : MUX2_X1 port map( A => REGISTERS_1_2_port, B => n5872, S => n87, Z 
                           => n4378);
   U4147 : MUX2_X1 port map( A => REGISTERS_1_1_port, B => n5873, S => n87, Z 
                           => n4377);
   U4148 : MUX2_X1 port map( A => REGISTERS_1_0_port, B => n5874, S => n87, Z 
                           => n4376);
   U4149 : OAI21_X1 port map( B1 => n5875, B2 => n5878, A => n5744, ZN => n5877
                           );
   U4150 : MUX2_X1 port map( A => REGISTERS_2_63_port, B => n5810, S => n89, Z 
                           => n4375);
   U4151 : MUX2_X1 port map( A => REGISTERS_2_62_port, B => n5812, S => n89, Z 
                           => n4374);
   U4152 : MUX2_X1 port map( A => REGISTERS_2_61_port, B => n5813, S => n89, Z 
                           => n4373);
   U4153 : MUX2_X1 port map( A => REGISTERS_2_60_port, B => n5814, S => n89, Z 
                           => n4372);
   U4154 : MUX2_X1 port map( A => REGISTERS_2_59_port, B => n5815, S => n89, Z 
                           => n4371);
   U4155 : MUX2_X1 port map( A => REGISTERS_2_58_port, B => n5816, S => n89, Z 
                           => n4370);
   U4156 : MUX2_X1 port map( A => REGISTERS_2_57_port, B => n5817, S => n89, Z 
                           => n4369);
   U4157 : MUX2_X1 port map( A => REGISTERS_2_56_port, B => n5818, S => n89, Z 
                           => n4368);
   U4158 : MUX2_X1 port map( A => REGISTERS_2_55_port, B => n5819, S => n89, Z 
                           => n4367);
   U4159 : MUX2_X1 port map( A => REGISTERS_2_54_port, B => n5820, S => n89, Z 
                           => n4366);
   U4160 : MUX2_X1 port map( A => REGISTERS_2_53_port, B => n5821, S => n89, Z 
                           => n4365);
   U4161 : MUX2_X1 port map( A => REGISTERS_2_52_port, B => n5822, S => n89, Z 
                           => n4364);
   U4162 : MUX2_X1 port map( A => REGISTERS_2_51_port, B => n5823, S => n89, Z 
                           => n4363);
   U4163 : MUX2_X1 port map( A => REGISTERS_2_50_port, B => n5824, S => n89, Z 
                           => n4362);
   U4164 : MUX2_X1 port map( A => REGISTERS_2_49_port, B => n5825, S => n89, Z 
                           => n4361);
   U4165 : MUX2_X1 port map( A => REGISTERS_2_48_port, B => n5826, S => n89, Z 
                           => n4360);
   U4166 : MUX2_X1 port map( A => REGISTERS_2_47_port, B => n5827, S => n89, Z 
                           => n4359);
   U4167 : MUX2_X1 port map( A => REGISTERS_2_46_port, B => n5828, S => n89, Z 
                           => n4358);
   U4168 : MUX2_X1 port map( A => REGISTERS_2_45_port, B => n5829, S => n89, Z 
                           => n4357);
   U4169 : MUX2_X1 port map( A => REGISTERS_2_44_port, B => n5830, S => n89, Z 
                           => n4356);
   U4170 : MUX2_X1 port map( A => REGISTERS_2_43_port, B => n5831, S => n89, Z 
                           => n4355);
   U4171 : MUX2_X1 port map( A => REGISTERS_2_42_port, B => n5832, S => n89, Z 
                           => n4354);
   U4172 : MUX2_X1 port map( A => REGISTERS_2_41_port, B => n5833, S => n89, Z 
                           => n4353);
   U4173 : MUX2_X1 port map( A => REGISTERS_2_40_port, B => n5834, S => n89, Z 
                           => n4352);
   U4174 : MUX2_X1 port map( A => REGISTERS_2_39_port, B => n5835, S => n89, Z 
                           => n4351);
   U4175 : MUX2_X1 port map( A => REGISTERS_2_38_port, B => n5836, S => n89, Z 
                           => n4350);
   U4176 : MUX2_X1 port map( A => REGISTERS_2_37_port, B => n5837, S => n89, Z 
                           => n4349);
   U4177 : MUX2_X1 port map( A => REGISTERS_2_36_port, B => n5838, S => n89, Z 
                           => n4348);
   U4178 : MUX2_X1 port map( A => REGISTERS_2_35_port, B => n5839, S => n89, Z 
                           => n4347);
   U4179 : MUX2_X1 port map( A => REGISTERS_2_34_port, B => n5840, S => n89, Z 
                           => n4346);
   U4180 : MUX2_X1 port map( A => REGISTERS_2_33_port, B => n5841, S => n89, Z 
                           => n4345);
   U4181 : MUX2_X1 port map( A => REGISTERS_2_32_port, B => n5842, S => n89, Z 
                           => n4344);
   U4182 : MUX2_X1 port map( A => REGISTERS_2_31_port, B => n5843, S => n89, Z 
                           => n4343);
   U4183 : MUX2_X1 port map( A => REGISTERS_2_30_port, B => n5844, S => n89, Z 
                           => n4342);
   U4184 : MUX2_X1 port map( A => REGISTERS_2_29_port, B => n5845, S => n89, Z 
                           => n4341);
   U4185 : MUX2_X1 port map( A => REGISTERS_2_28_port, B => n5846, S => n89, Z 
                           => n4340);
   U4186 : MUX2_X1 port map( A => REGISTERS_2_27_port, B => n5847, S => n89, Z 
                           => n4339);
   U4187 : MUX2_X1 port map( A => REGISTERS_2_26_port, B => n5848, S => n89, Z 
                           => n4338);
   U4188 : MUX2_X1 port map( A => REGISTERS_2_25_port, B => n5849, S => n89, Z 
                           => n4337);
   U4189 : MUX2_X1 port map( A => REGISTERS_2_24_port, B => n5850, S => n89, Z 
                           => n4336);
   U4190 : MUX2_X1 port map( A => REGISTERS_2_23_port, B => n5851, S => n89, Z 
                           => n4335);
   U4191 : MUX2_X1 port map( A => REGISTERS_2_22_port, B => n5852, S => n89, Z 
                           => n4334);
   U4192 : MUX2_X1 port map( A => REGISTERS_2_21_port, B => n5853, S => n89, Z 
                           => n4333);
   U4193 : MUX2_X1 port map( A => REGISTERS_2_20_port, B => n5854, S => n89, Z 
                           => n4332);
   U4194 : MUX2_X1 port map( A => REGISTERS_2_19_port, B => n5855, S => n89, Z 
                           => n4331);
   U4195 : MUX2_X1 port map( A => REGISTERS_2_18_port, B => n5856, S => n89, Z 
                           => n4330);
   U4196 : MUX2_X1 port map( A => REGISTERS_2_17_port, B => n5857, S => n89, Z 
                           => n4329);
   U4197 : MUX2_X1 port map( A => REGISTERS_2_16_port, B => n5858, S => n89, Z 
                           => n4328);
   U4198 : MUX2_X1 port map( A => REGISTERS_2_15_port, B => n5859, S => n89, Z 
                           => n4327);
   U4199 : MUX2_X1 port map( A => REGISTERS_2_14_port, B => n5860, S => n89, Z 
                           => n4326);
   U4200 : MUX2_X1 port map( A => REGISTERS_2_13_port, B => n5861, S => n89, Z 
                           => n4325);
   U4201 : MUX2_X1 port map( A => REGISTERS_2_12_port, B => n5862, S => n89, Z 
                           => n4324);
   U4202 : MUX2_X1 port map( A => REGISTERS_2_11_port, B => n5863, S => n89, Z 
                           => n4323);
   U4203 : MUX2_X1 port map( A => REGISTERS_2_10_port, B => n5864, S => n89, Z 
                           => n4322);
   U4204 : MUX2_X1 port map( A => REGISTERS_2_9_port, B => n5865, S => n89, Z 
                           => n4321);
   U4205 : MUX2_X1 port map( A => REGISTERS_2_8_port, B => n5866, S => n89, Z 
                           => n4320);
   U4206 : MUX2_X1 port map( A => REGISTERS_2_7_port, B => n5867, S => n89, Z 
                           => n4319);
   U4207 : MUX2_X1 port map( A => REGISTERS_2_6_port, B => n5868, S => n89, Z 
                           => n4318);
   U4208 : MUX2_X1 port map( A => REGISTERS_2_5_port, B => n5869, S => n89, Z 
                           => n4317);
   U4209 : MUX2_X1 port map( A => REGISTERS_2_4_port, B => n5870, S => n89, Z 
                           => n4316);
   U4210 : MUX2_X1 port map( A => REGISTERS_2_3_port, B => n5871, S => n89, Z 
                           => n4315);
   U4211 : MUX2_X1 port map( A => REGISTERS_2_2_port, B => n5872, S => n89, Z 
                           => n4314);
   U4212 : MUX2_X1 port map( A => REGISTERS_2_1_port, B => n5873, S => n89, Z 
                           => n4313);
   U4213 : MUX2_X1 port map( A => REGISTERS_2_0_port, B => n5874, S => n89, Z 
                           => n4312);
   U4214 : OAI21_X1 port map( B1 => n5875, B2 => n5880, A => n5744, ZN => n5879
                           );
   U4215 : MUX2_X1 port map( A => REGISTERS_3_63_port, B => n5810, S => n77, Z 
                           => n4311);
   U4216 : MUX2_X1 port map( A => REGISTERS_3_62_port, B => n5812, S => n77, Z 
                           => n4310);
   U4217 : MUX2_X1 port map( A => REGISTERS_3_61_port, B => n5813, S => n77, Z 
                           => n4309);
   U4218 : MUX2_X1 port map( A => REGISTERS_3_60_port, B => n5814, S => n77, Z 
                           => n4308);
   U4219 : MUX2_X1 port map( A => REGISTERS_3_59_port, B => n5815, S => n77, Z 
                           => n4307);
   U4220 : MUX2_X1 port map( A => REGISTERS_3_58_port, B => n5816, S => n77, Z 
                           => n4306);
   U4221 : MUX2_X1 port map( A => REGISTERS_3_57_port, B => n5817, S => n77, Z 
                           => n4305);
   U4222 : MUX2_X1 port map( A => REGISTERS_3_56_port, B => n5818, S => n77, Z 
                           => n4304);
   U4223 : MUX2_X1 port map( A => REGISTERS_3_55_port, B => n5819, S => n77, Z 
                           => n4303);
   U4224 : MUX2_X1 port map( A => REGISTERS_3_54_port, B => n5820, S => n77, Z 
                           => n4302);
   U4225 : MUX2_X1 port map( A => REGISTERS_3_53_port, B => n5821, S => n77, Z 
                           => n4301);
   U4226 : MUX2_X1 port map( A => REGISTERS_3_52_port, B => n5822, S => n77, Z 
                           => n4300);
   U4227 : MUX2_X1 port map( A => REGISTERS_3_51_port, B => n5823, S => n77, Z 
                           => n4299);
   U4228 : MUX2_X1 port map( A => REGISTERS_3_50_port, B => n5824, S => n77, Z 
                           => n4298);
   U4229 : MUX2_X1 port map( A => REGISTERS_3_49_port, B => n5825, S => n77, Z 
                           => n4297);
   U4230 : MUX2_X1 port map( A => REGISTERS_3_48_port, B => n5826, S => n77, Z 
                           => n4296);
   U4231 : MUX2_X1 port map( A => REGISTERS_3_47_port, B => n5827, S => n77, Z 
                           => n4295);
   U4232 : MUX2_X1 port map( A => REGISTERS_3_46_port, B => n5828, S => n77, Z 
                           => n4294);
   U4233 : MUX2_X1 port map( A => REGISTERS_3_45_port, B => n5829, S => n77, Z 
                           => n4293);
   U4234 : MUX2_X1 port map( A => REGISTERS_3_44_port, B => n5830, S => n77, Z 
                           => n4292);
   U4235 : MUX2_X1 port map( A => REGISTERS_3_43_port, B => n5831, S => n77, Z 
                           => n4291);
   U4236 : MUX2_X1 port map( A => REGISTERS_3_42_port, B => n5832, S => n77, Z 
                           => n4290);
   U4237 : MUX2_X1 port map( A => REGISTERS_3_41_port, B => n5833, S => n77, Z 
                           => n4289);
   U4238 : MUX2_X1 port map( A => REGISTERS_3_40_port, B => n5834, S => n77, Z 
                           => n4288);
   U4239 : MUX2_X1 port map( A => REGISTERS_3_39_port, B => n5835, S => n77, Z 
                           => n4287);
   U4240 : MUX2_X1 port map( A => REGISTERS_3_38_port, B => n5836, S => n77, Z 
                           => n4286);
   U4241 : MUX2_X1 port map( A => REGISTERS_3_37_port, B => n5837, S => n77, Z 
                           => n4285);
   U4242 : MUX2_X1 port map( A => REGISTERS_3_36_port, B => n5838, S => n77, Z 
                           => n4284);
   U4243 : MUX2_X1 port map( A => REGISTERS_3_35_port, B => n5839, S => n77, Z 
                           => n4283);
   U4244 : MUX2_X1 port map( A => REGISTERS_3_34_port, B => n5840, S => n77, Z 
                           => n4282);
   U4245 : MUX2_X1 port map( A => REGISTERS_3_33_port, B => n5841, S => n77, Z 
                           => n4281);
   U4246 : MUX2_X1 port map( A => REGISTERS_3_32_port, B => n5842, S => n77, Z 
                           => n4280);
   U4247 : MUX2_X1 port map( A => REGISTERS_3_31_port, B => n5843, S => n77, Z 
                           => n4279);
   U4248 : MUX2_X1 port map( A => REGISTERS_3_30_port, B => n5844, S => n77, Z 
                           => n4278);
   U4249 : MUX2_X1 port map( A => REGISTERS_3_29_port, B => n5845, S => n77, Z 
                           => n4277);
   U4250 : MUX2_X1 port map( A => REGISTERS_3_28_port, B => n5846, S => n77, Z 
                           => n4276);
   U4251 : MUX2_X1 port map( A => REGISTERS_3_27_port, B => n5847, S => n77, Z 
                           => n4275);
   U4252 : MUX2_X1 port map( A => REGISTERS_3_26_port, B => n5848, S => n77, Z 
                           => n4274);
   U4253 : MUX2_X1 port map( A => REGISTERS_3_25_port, B => n5849, S => n77, Z 
                           => n4273);
   U4254 : MUX2_X1 port map( A => REGISTERS_3_24_port, B => n5850, S => n77, Z 
                           => n4272);
   U4255 : MUX2_X1 port map( A => REGISTERS_3_23_port, B => n5851, S => n77, Z 
                           => n4271);
   U4256 : MUX2_X1 port map( A => REGISTERS_3_22_port, B => n5852, S => n77, Z 
                           => n4270);
   U4257 : MUX2_X1 port map( A => REGISTERS_3_21_port, B => n5853, S => n77, Z 
                           => n4269);
   U4258 : MUX2_X1 port map( A => REGISTERS_3_20_port, B => n5854, S => n77, Z 
                           => n4268);
   U4259 : MUX2_X1 port map( A => REGISTERS_3_19_port, B => n5855, S => n77, Z 
                           => n4267);
   U4260 : MUX2_X1 port map( A => REGISTERS_3_18_port, B => n5856, S => n77, Z 
                           => n4266);
   U4261 : MUX2_X1 port map( A => REGISTERS_3_17_port, B => n5857, S => n77, Z 
                           => n4265);
   U4262 : MUX2_X1 port map( A => REGISTERS_3_16_port, B => n5858, S => n77, Z 
                           => n4264);
   U4263 : MUX2_X1 port map( A => REGISTERS_3_15_port, B => n5859, S => n77, Z 
                           => n4263);
   U4264 : MUX2_X1 port map( A => REGISTERS_3_14_port, B => n5860, S => n77, Z 
                           => n4262);
   U4265 : MUX2_X1 port map( A => REGISTERS_3_13_port, B => n5861, S => n77, Z 
                           => n4261);
   U4266 : MUX2_X1 port map( A => REGISTERS_3_12_port, B => n5862, S => n77, Z 
                           => n4260);
   U4267 : MUX2_X1 port map( A => REGISTERS_3_11_port, B => n5863, S => n77, Z 
                           => n4259);
   U4268 : MUX2_X1 port map( A => REGISTERS_3_10_port, B => n5864, S => n77, Z 
                           => n4258);
   U4269 : MUX2_X1 port map( A => REGISTERS_3_9_port, B => n5865, S => n77, Z 
                           => n4257);
   U4270 : MUX2_X1 port map( A => REGISTERS_3_8_port, B => n5866, S => n77, Z 
                           => n4256);
   U4271 : MUX2_X1 port map( A => REGISTERS_3_7_port, B => n5867, S => n77, Z 
                           => n4255);
   U4272 : MUX2_X1 port map( A => REGISTERS_3_6_port, B => n5868, S => n77, Z 
                           => n4254);
   U4273 : MUX2_X1 port map( A => REGISTERS_3_5_port, B => n5869, S => n77, Z 
                           => n4253);
   U4274 : MUX2_X1 port map( A => REGISTERS_3_4_port, B => n5870, S => n77, Z 
                           => n4252);
   U4275 : MUX2_X1 port map( A => REGISTERS_3_3_port, B => n5871, S => n77, Z 
                           => n4251);
   U4276 : MUX2_X1 port map( A => REGISTERS_3_2_port, B => n5872, S => n77, Z 
                           => n4250);
   U4277 : MUX2_X1 port map( A => REGISTERS_3_1_port, B => n5873, S => n77, Z 
                           => n4249);
   U4278 : MUX2_X1 port map( A => REGISTERS_3_0_port, B => n5874, S => n77, Z 
                           => n4248);
   U4279 : OAI21_X1 port map( B1 => n5875, B2 => n5882, A => n5744, ZN => n5881
                           );
   U4280 : MUX2_X1 port map( A => REGISTERS_4_63_port, B => n5810, S => n79, Z 
                           => n4247);
   U4281 : MUX2_X1 port map( A => REGISTERS_4_62_port, B => n5812, S => n79, Z 
                           => n4246);
   U4282 : MUX2_X1 port map( A => REGISTERS_4_61_port, B => n5813, S => n79, Z 
                           => n4245);
   U4283 : MUX2_X1 port map( A => REGISTERS_4_60_port, B => n5814, S => n79, Z 
                           => n4244);
   U4284 : MUX2_X1 port map( A => REGISTERS_4_59_port, B => n5815, S => n79, Z 
                           => n4243);
   U4285 : MUX2_X1 port map( A => REGISTERS_4_58_port, B => n5816, S => n79, Z 
                           => n4242);
   U4286 : MUX2_X1 port map( A => REGISTERS_4_57_port, B => n5817, S => n79, Z 
                           => n4241);
   U4287 : MUX2_X1 port map( A => REGISTERS_4_56_port, B => n5818, S => n79, Z 
                           => n4240);
   U4288 : MUX2_X1 port map( A => REGISTERS_4_55_port, B => n5819, S => n79, Z 
                           => n4239);
   U4289 : MUX2_X1 port map( A => REGISTERS_4_54_port, B => n5820, S => n79, Z 
                           => n4238);
   U4290 : MUX2_X1 port map( A => REGISTERS_4_53_port, B => n5821, S => n79, Z 
                           => n4237);
   U4291 : MUX2_X1 port map( A => REGISTERS_4_52_port, B => n5822, S => n79, Z 
                           => n4236);
   U4292 : MUX2_X1 port map( A => REGISTERS_4_51_port, B => n5823, S => n79, Z 
                           => n4235);
   U4293 : MUX2_X1 port map( A => REGISTERS_4_50_port, B => n5824, S => n79, Z 
                           => n4234);
   U4294 : MUX2_X1 port map( A => REGISTERS_4_49_port, B => n5825, S => n79, Z 
                           => n4233);
   U4295 : MUX2_X1 port map( A => REGISTERS_4_48_port, B => n5826, S => n79, Z 
                           => n4232);
   U4296 : MUX2_X1 port map( A => REGISTERS_4_47_port, B => n5827, S => n79, Z 
                           => n4231);
   U4297 : MUX2_X1 port map( A => REGISTERS_4_46_port, B => n5828, S => n79, Z 
                           => n4230);
   U4298 : MUX2_X1 port map( A => REGISTERS_4_45_port, B => n5829, S => n79, Z 
                           => n4229);
   U4299 : MUX2_X1 port map( A => REGISTERS_4_44_port, B => n5830, S => n79, Z 
                           => n4228);
   U4300 : MUX2_X1 port map( A => REGISTERS_4_43_port, B => n5831, S => n79, Z 
                           => n4227);
   U4301 : MUX2_X1 port map( A => REGISTERS_4_42_port, B => n5832, S => n79, Z 
                           => n4226);
   U4302 : MUX2_X1 port map( A => REGISTERS_4_41_port, B => n5833, S => n79, Z 
                           => n4225);
   U4303 : MUX2_X1 port map( A => REGISTERS_4_40_port, B => n5834, S => n79, Z 
                           => n4224);
   U4304 : MUX2_X1 port map( A => REGISTERS_4_39_port, B => n5835, S => n79, Z 
                           => n4223);
   U4305 : MUX2_X1 port map( A => REGISTERS_4_38_port, B => n5836, S => n79, Z 
                           => n4222);
   U4306 : MUX2_X1 port map( A => REGISTERS_4_37_port, B => n5837, S => n79, Z 
                           => n4221);
   U4307 : MUX2_X1 port map( A => REGISTERS_4_36_port, B => n5838, S => n79, Z 
                           => n4220);
   U4308 : MUX2_X1 port map( A => REGISTERS_4_35_port, B => n5839, S => n79, Z 
                           => n4219);
   U4309 : MUX2_X1 port map( A => REGISTERS_4_34_port, B => n5840, S => n79, Z 
                           => n4218);
   U4310 : MUX2_X1 port map( A => REGISTERS_4_33_port, B => n5841, S => n79, Z 
                           => n4217);
   U4311 : MUX2_X1 port map( A => REGISTERS_4_32_port, B => n5842, S => n79, Z 
                           => n4216);
   U4312 : MUX2_X1 port map( A => REGISTERS_4_31_port, B => n5843, S => n79, Z 
                           => n4215);
   U4313 : MUX2_X1 port map( A => REGISTERS_4_30_port, B => n5844, S => n79, Z 
                           => n4214);
   U4314 : MUX2_X1 port map( A => REGISTERS_4_29_port, B => n5845, S => n79, Z 
                           => n4213);
   U4315 : MUX2_X1 port map( A => REGISTERS_4_28_port, B => n5846, S => n79, Z 
                           => n4212);
   U4316 : MUX2_X1 port map( A => REGISTERS_4_27_port, B => n5847, S => n79, Z 
                           => n4211);
   U4317 : MUX2_X1 port map( A => REGISTERS_4_26_port, B => n5848, S => n79, Z 
                           => n4210);
   U4318 : MUX2_X1 port map( A => REGISTERS_4_25_port, B => n5849, S => n79, Z 
                           => n4209);
   U4319 : MUX2_X1 port map( A => REGISTERS_4_24_port, B => n5850, S => n79, Z 
                           => n4208);
   U4320 : MUX2_X1 port map( A => REGISTERS_4_23_port, B => n5851, S => n79, Z 
                           => n4207);
   U4321 : MUX2_X1 port map( A => REGISTERS_4_22_port, B => n5852, S => n79, Z 
                           => n4206);
   U4322 : MUX2_X1 port map( A => REGISTERS_4_21_port, B => n5853, S => n79, Z 
                           => n4205);
   U4323 : MUX2_X1 port map( A => REGISTERS_4_20_port, B => n5854, S => n79, Z 
                           => n4204);
   U4324 : MUX2_X1 port map( A => REGISTERS_4_19_port, B => n5855, S => n79, Z 
                           => n4203);
   U4325 : MUX2_X1 port map( A => REGISTERS_4_18_port, B => n5856, S => n79, Z 
                           => n4202);
   U4326 : MUX2_X1 port map( A => REGISTERS_4_17_port, B => n5857, S => n79, Z 
                           => n4201);
   U4327 : MUX2_X1 port map( A => REGISTERS_4_16_port, B => n5858, S => n79, Z 
                           => n4200);
   U4328 : MUX2_X1 port map( A => REGISTERS_4_15_port, B => n5859, S => n79, Z 
                           => n4199);
   U4329 : MUX2_X1 port map( A => REGISTERS_4_14_port, B => n5860, S => n79, Z 
                           => n4198);
   U4330 : MUX2_X1 port map( A => REGISTERS_4_13_port, B => n5861, S => n79, Z 
                           => n4197);
   U4331 : MUX2_X1 port map( A => REGISTERS_4_12_port, B => n5862, S => n79, Z 
                           => n4196);
   U4332 : MUX2_X1 port map( A => REGISTERS_4_11_port, B => n5863, S => n79, Z 
                           => n4195);
   U4333 : MUX2_X1 port map( A => REGISTERS_4_10_port, B => n5864, S => n79, Z 
                           => n4194);
   U4334 : MUX2_X1 port map( A => REGISTERS_4_9_port, B => n5865, S => n79, Z 
                           => n4193);
   U4335 : MUX2_X1 port map( A => REGISTERS_4_8_port, B => n5866, S => n79, Z 
                           => n4192);
   U4336 : MUX2_X1 port map( A => REGISTERS_4_7_port, B => n5867, S => n79, Z 
                           => n4191);
   U4337 : MUX2_X1 port map( A => REGISTERS_4_6_port, B => n5868, S => n79, Z 
                           => n4190);
   U4338 : MUX2_X1 port map( A => REGISTERS_4_5_port, B => n5869, S => n79, Z 
                           => n4189);
   U4339 : MUX2_X1 port map( A => REGISTERS_4_4_port, B => n5870, S => n79, Z 
                           => n4188);
   U4340 : MUX2_X1 port map( A => REGISTERS_4_3_port, B => n5871, S => n79, Z 
                           => n4187);
   U4341 : MUX2_X1 port map( A => REGISTERS_4_2_port, B => n5872, S => n79, Z 
                           => n4186);
   U4342 : MUX2_X1 port map( A => REGISTERS_4_1_port, B => n5873, S => n79, Z 
                           => n4185);
   U4343 : MUX2_X1 port map( A => REGISTERS_4_0_port, B => n5874, S => n79, Z 
                           => n4184);
   U4344 : OAI21_X1 port map( B1 => n5875, B2 => n5884, A => n5744, ZN => n5883
                           );
   U4345 : MUX2_X1 port map( A => REGISTERS_5_63_port, B => n5810, S => n81, Z 
                           => n4183);
   U4346 : MUX2_X1 port map( A => REGISTERS_5_62_port, B => n5812, S => n81, Z 
                           => n4182);
   U4347 : MUX2_X1 port map( A => REGISTERS_5_61_port, B => n5813, S => n81, Z 
                           => n4181);
   U4348 : MUX2_X1 port map( A => REGISTERS_5_60_port, B => n5814, S => n81, Z 
                           => n4180);
   U4349 : MUX2_X1 port map( A => REGISTERS_5_59_port, B => n5815, S => n81, Z 
                           => n4179);
   U4350 : MUX2_X1 port map( A => REGISTERS_5_58_port, B => n5816, S => n81, Z 
                           => n4178);
   U4351 : MUX2_X1 port map( A => REGISTERS_5_57_port, B => n5817, S => n81, Z 
                           => n4177);
   U4352 : MUX2_X1 port map( A => REGISTERS_5_56_port, B => n5818, S => n81, Z 
                           => n4176);
   U4353 : MUX2_X1 port map( A => REGISTERS_5_55_port, B => n5819, S => n81, Z 
                           => n4175);
   U4354 : MUX2_X1 port map( A => REGISTERS_5_54_port, B => n5820, S => n81, Z 
                           => n4174);
   U4355 : MUX2_X1 port map( A => REGISTERS_5_53_port, B => n5821, S => n81, Z 
                           => n4173);
   U4356 : MUX2_X1 port map( A => REGISTERS_5_52_port, B => n5822, S => n81, Z 
                           => n4172);
   U4357 : MUX2_X1 port map( A => REGISTERS_5_51_port, B => n5823, S => n81, Z 
                           => n4171);
   U4358 : MUX2_X1 port map( A => REGISTERS_5_50_port, B => n5824, S => n81, Z 
                           => n4170);
   U4359 : MUX2_X1 port map( A => REGISTERS_5_49_port, B => n5825, S => n81, Z 
                           => n4169);
   U4360 : MUX2_X1 port map( A => REGISTERS_5_48_port, B => n5826, S => n81, Z 
                           => n4168);
   U4361 : MUX2_X1 port map( A => REGISTERS_5_47_port, B => n5827, S => n81, Z 
                           => n4167);
   U4362 : MUX2_X1 port map( A => REGISTERS_5_46_port, B => n5828, S => n81, Z 
                           => n4166);
   U4363 : MUX2_X1 port map( A => REGISTERS_5_45_port, B => n5829, S => n81, Z 
                           => n4165);
   U4364 : MUX2_X1 port map( A => REGISTERS_5_44_port, B => n5830, S => n81, Z 
                           => n4164);
   U4365 : MUX2_X1 port map( A => REGISTERS_5_43_port, B => n5831, S => n81, Z 
                           => n4163);
   U4366 : MUX2_X1 port map( A => REGISTERS_5_42_port, B => n5832, S => n81, Z 
                           => n4162);
   U4367 : MUX2_X1 port map( A => REGISTERS_5_41_port, B => n5833, S => n81, Z 
                           => n4161);
   U4368 : MUX2_X1 port map( A => REGISTERS_5_40_port, B => n5834, S => n81, Z 
                           => n4160);
   U4369 : MUX2_X1 port map( A => REGISTERS_5_39_port, B => n5835, S => n81, Z 
                           => n4159);
   U4370 : MUX2_X1 port map( A => REGISTERS_5_38_port, B => n5836, S => n81, Z 
                           => n4158);
   U4371 : MUX2_X1 port map( A => REGISTERS_5_37_port, B => n5837, S => n81, Z 
                           => n4157);
   U4372 : MUX2_X1 port map( A => REGISTERS_5_36_port, B => n5838, S => n81, Z 
                           => n4156);
   U4373 : MUX2_X1 port map( A => REGISTERS_5_35_port, B => n5839, S => n81, Z 
                           => n4155);
   U4374 : MUX2_X1 port map( A => REGISTERS_5_34_port, B => n5840, S => n81, Z 
                           => n4154);
   U4375 : MUX2_X1 port map( A => REGISTERS_5_33_port, B => n5841, S => n81, Z 
                           => n4153);
   U4376 : MUX2_X1 port map( A => REGISTERS_5_32_port, B => n5842, S => n81, Z 
                           => n4152);
   U4377 : MUX2_X1 port map( A => REGISTERS_5_31_port, B => n5843, S => n81, Z 
                           => n4151);
   U4378 : MUX2_X1 port map( A => REGISTERS_5_30_port, B => n5844, S => n81, Z 
                           => n4150);
   U4379 : MUX2_X1 port map( A => REGISTERS_5_29_port, B => n5845, S => n81, Z 
                           => n4149);
   U4380 : MUX2_X1 port map( A => REGISTERS_5_28_port, B => n5846, S => n81, Z 
                           => n4148);
   U4381 : MUX2_X1 port map( A => REGISTERS_5_27_port, B => n5847, S => n81, Z 
                           => n4147);
   U4382 : MUX2_X1 port map( A => REGISTERS_5_26_port, B => n5848, S => n81, Z 
                           => n4146);
   U4383 : MUX2_X1 port map( A => REGISTERS_5_25_port, B => n5849, S => n81, Z 
                           => n4145);
   U4384 : MUX2_X1 port map( A => REGISTERS_5_24_port, B => n5850, S => n81, Z 
                           => n4144);
   U4385 : MUX2_X1 port map( A => REGISTERS_5_23_port, B => n5851, S => n81, Z 
                           => n4143);
   U4386 : MUX2_X1 port map( A => REGISTERS_5_22_port, B => n5852, S => n81, Z 
                           => n4142);
   U4387 : MUX2_X1 port map( A => REGISTERS_5_21_port, B => n5853, S => n81, Z 
                           => n4141);
   U4388 : MUX2_X1 port map( A => REGISTERS_5_20_port, B => n5854, S => n81, Z 
                           => n4140);
   U4389 : MUX2_X1 port map( A => REGISTERS_5_19_port, B => n5855, S => n81, Z 
                           => n4139);
   U4390 : MUX2_X1 port map( A => REGISTERS_5_18_port, B => n5856, S => n81, Z 
                           => n4138);
   U4391 : MUX2_X1 port map( A => REGISTERS_5_17_port, B => n5857, S => n81, Z 
                           => n4137);
   U4392 : MUX2_X1 port map( A => REGISTERS_5_16_port, B => n5858, S => n81, Z 
                           => n4136);
   U4393 : MUX2_X1 port map( A => REGISTERS_5_15_port, B => n5859, S => n81, Z 
                           => n4135);
   U4394 : MUX2_X1 port map( A => REGISTERS_5_14_port, B => n5860, S => n81, Z 
                           => n4134);
   U4395 : MUX2_X1 port map( A => REGISTERS_5_13_port, B => n5861, S => n81, Z 
                           => n4133);
   U4396 : MUX2_X1 port map( A => REGISTERS_5_12_port, B => n5862, S => n81, Z 
                           => n4132);
   U4397 : MUX2_X1 port map( A => REGISTERS_5_11_port, B => n5863, S => n81, Z 
                           => n4131);
   U4398 : MUX2_X1 port map( A => REGISTERS_5_10_port, B => n5864, S => n81, Z 
                           => n4130);
   U4399 : MUX2_X1 port map( A => REGISTERS_5_9_port, B => n5865, S => n81, Z 
                           => n4129);
   U4400 : MUX2_X1 port map( A => REGISTERS_5_8_port, B => n5866, S => n81, Z 
                           => n4128);
   U4401 : MUX2_X1 port map( A => REGISTERS_5_7_port, B => n5867, S => n81, Z 
                           => n4127);
   U4402 : MUX2_X1 port map( A => REGISTERS_5_6_port, B => n5868, S => n81, Z 
                           => n4126);
   U4403 : MUX2_X1 port map( A => REGISTERS_5_5_port, B => n5869, S => n81, Z 
                           => n4125);
   U4404 : MUX2_X1 port map( A => REGISTERS_5_4_port, B => n5870, S => n81, Z 
                           => n4124);
   U4405 : MUX2_X1 port map( A => REGISTERS_5_3_port, B => n5871, S => n81, Z 
                           => n4123);
   U4406 : MUX2_X1 port map( A => REGISTERS_5_2_port, B => n5872, S => n81, Z 
                           => n4122);
   U4407 : MUX2_X1 port map( A => REGISTERS_5_1_port, B => n5873, S => n81, Z 
                           => n4121);
   U4408 : MUX2_X1 port map( A => REGISTERS_5_0_port, B => n5874, S => n81, Z 
                           => n4120);
   U4409 : OAI21_X1 port map( B1 => n5875, B2 => n5886, A => n5744, ZN => n5885
                           );
   U4410 : MUX2_X1 port map( A => REGISTERS_6_63_port, B => n5810, S => n83, Z 
                           => n4119);
   U4411 : MUX2_X1 port map( A => REGISTERS_6_62_port, B => n5812, S => n83, Z 
                           => n4118);
   U4412 : MUX2_X1 port map( A => REGISTERS_6_61_port, B => n5813, S => n83, Z 
                           => n4117);
   U4413 : MUX2_X1 port map( A => REGISTERS_6_60_port, B => n5814, S => n83, Z 
                           => n4116);
   U4414 : MUX2_X1 port map( A => REGISTERS_6_59_port, B => n5815, S => n83, Z 
                           => n4115);
   U4415 : MUX2_X1 port map( A => REGISTERS_6_58_port, B => n5816, S => n83, Z 
                           => n4114);
   U4416 : MUX2_X1 port map( A => REGISTERS_6_57_port, B => n5817, S => n83, Z 
                           => n4113);
   U4417 : MUX2_X1 port map( A => REGISTERS_6_56_port, B => n5818, S => n83, Z 
                           => n4112);
   U4418 : MUX2_X1 port map( A => REGISTERS_6_55_port, B => n5819, S => n83, Z 
                           => n4111);
   U4419 : MUX2_X1 port map( A => REGISTERS_6_54_port, B => n5820, S => n83, Z 
                           => n4110);
   U4420 : MUX2_X1 port map( A => REGISTERS_6_53_port, B => n5821, S => n83, Z 
                           => n4109);
   U4421 : MUX2_X1 port map( A => REGISTERS_6_52_port, B => n5822, S => n83, Z 
                           => n4108);
   U4422 : MUX2_X1 port map( A => REGISTERS_6_51_port, B => n5823, S => n83, Z 
                           => n4107);
   U4423 : MUX2_X1 port map( A => REGISTERS_6_50_port, B => n5824, S => n83, Z 
                           => n4106);
   U4424 : MUX2_X1 port map( A => REGISTERS_6_49_port, B => n5825, S => n83, Z 
                           => n4105);
   U4425 : MUX2_X1 port map( A => REGISTERS_6_48_port, B => n5826, S => n83, Z 
                           => n4104);
   U4426 : MUX2_X1 port map( A => REGISTERS_6_47_port, B => n5827, S => n83, Z 
                           => n4103);
   U4427 : MUX2_X1 port map( A => REGISTERS_6_46_port, B => n5828, S => n83, Z 
                           => n4102);
   U4428 : MUX2_X1 port map( A => REGISTERS_6_45_port, B => n5829, S => n83, Z 
                           => n4101);
   U4429 : MUX2_X1 port map( A => REGISTERS_6_44_port, B => n5830, S => n83, Z 
                           => n4100);
   U4430 : MUX2_X1 port map( A => REGISTERS_6_43_port, B => n5831, S => n83, Z 
                           => n4099);
   U4431 : MUX2_X1 port map( A => REGISTERS_6_42_port, B => n5832, S => n83, Z 
                           => n4098);
   U4432 : MUX2_X1 port map( A => REGISTERS_6_41_port, B => n5833, S => n83, Z 
                           => n4097);
   U4433 : MUX2_X1 port map( A => REGISTERS_6_40_port, B => n5834, S => n83, Z 
                           => n4096);
   U4434 : MUX2_X1 port map( A => REGISTERS_6_39_port, B => n5835, S => n83, Z 
                           => n4095);
   U4435 : MUX2_X1 port map( A => REGISTERS_6_38_port, B => n5836, S => n83, Z 
                           => n4094);
   U4436 : MUX2_X1 port map( A => REGISTERS_6_37_port, B => n5837, S => n83, Z 
                           => n4093);
   U4437 : MUX2_X1 port map( A => REGISTERS_6_36_port, B => n5838, S => n83, Z 
                           => n4092);
   U4438 : MUX2_X1 port map( A => REGISTERS_6_35_port, B => n5839, S => n83, Z 
                           => n4091);
   U4439 : MUX2_X1 port map( A => REGISTERS_6_34_port, B => n5840, S => n83, Z 
                           => n4090);
   U4440 : MUX2_X1 port map( A => REGISTERS_6_33_port, B => n5841, S => n83, Z 
                           => n4089);
   U4441 : MUX2_X1 port map( A => REGISTERS_6_32_port, B => n5842, S => n83, Z 
                           => n4088);
   U4442 : MUX2_X1 port map( A => REGISTERS_6_31_port, B => n5843, S => n83, Z 
                           => n4087);
   U4443 : MUX2_X1 port map( A => REGISTERS_6_30_port, B => n5844, S => n83, Z 
                           => n4086);
   U4444 : MUX2_X1 port map( A => REGISTERS_6_29_port, B => n5845, S => n83, Z 
                           => n4085);
   U4445 : MUX2_X1 port map( A => REGISTERS_6_28_port, B => n5846, S => n83, Z 
                           => n4084);
   U4446 : MUX2_X1 port map( A => REGISTERS_6_27_port, B => n5847, S => n83, Z 
                           => n4083);
   U4447 : MUX2_X1 port map( A => REGISTERS_6_26_port, B => n5848, S => n83, Z 
                           => n4082);
   U4448 : MUX2_X1 port map( A => REGISTERS_6_25_port, B => n5849, S => n83, Z 
                           => n4081);
   U4449 : MUX2_X1 port map( A => REGISTERS_6_24_port, B => n5850, S => n83, Z 
                           => n4080);
   U4450 : MUX2_X1 port map( A => REGISTERS_6_23_port, B => n5851, S => n83, Z 
                           => n4079);
   U4451 : MUX2_X1 port map( A => REGISTERS_6_22_port, B => n5852, S => n83, Z 
                           => n4078);
   U4452 : MUX2_X1 port map( A => REGISTERS_6_21_port, B => n5853, S => n83, Z 
                           => n4077);
   U4453 : MUX2_X1 port map( A => REGISTERS_6_20_port, B => n5854, S => n83, Z 
                           => n4076);
   U4454 : MUX2_X1 port map( A => REGISTERS_6_19_port, B => n5855, S => n83, Z 
                           => n4075);
   U4455 : MUX2_X1 port map( A => REGISTERS_6_18_port, B => n5856, S => n83, Z 
                           => n4074);
   U4456 : MUX2_X1 port map( A => REGISTERS_6_17_port, B => n5857, S => n83, Z 
                           => n4073);
   U4457 : MUX2_X1 port map( A => REGISTERS_6_16_port, B => n5858, S => n83, Z 
                           => n4072);
   U4458 : MUX2_X1 port map( A => REGISTERS_6_15_port, B => n5859, S => n83, Z 
                           => n4071);
   U4459 : MUX2_X1 port map( A => REGISTERS_6_14_port, B => n5860, S => n83, Z 
                           => n4070);
   U4460 : MUX2_X1 port map( A => REGISTERS_6_13_port, B => n5861, S => n83, Z 
                           => n4069);
   U4461 : MUX2_X1 port map( A => REGISTERS_6_12_port, B => n5862, S => n83, Z 
                           => n4068);
   U4462 : MUX2_X1 port map( A => REGISTERS_6_11_port, B => n5863, S => n83, Z 
                           => n4067);
   U4463 : MUX2_X1 port map( A => REGISTERS_6_10_port, B => n5864, S => n83, Z 
                           => n4066);
   U4464 : MUX2_X1 port map( A => REGISTERS_6_9_port, B => n5865, S => n83, Z 
                           => n4065);
   U4465 : MUX2_X1 port map( A => REGISTERS_6_8_port, B => n5866, S => n83, Z 
                           => n4064);
   U4466 : MUX2_X1 port map( A => REGISTERS_6_7_port, B => n5867, S => n83, Z 
                           => n4063);
   U4467 : MUX2_X1 port map( A => REGISTERS_6_6_port, B => n5868, S => n83, Z 
                           => n4062);
   U4468 : MUX2_X1 port map( A => REGISTERS_6_5_port, B => n5869, S => n83, Z 
                           => n4061);
   U4469 : MUX2_X1 port map( A => REGISTERS_6_4_port, B => n5870, S => n83, Z 
                           => n4060);
   U4470 : MUX2_X1 port map( A => REGISTERS_6_3_port, B => n5871, S => n83, Z 
                           => n4059);
   U4471 : MUX2_X1 port map( A => REGISTERS_6_2_port, B => n5872, S => n83, Z 
                           => n4058);
   U4472 : MUX2_X1 port map( A => REGISTERS_6_1_port, B => n5873, S => n83, Z 
                           => n4057);
   U4473 : MUX2_X1 port map( A => REGISTERS_6_0_port, B => n5874, S => n83, Z 
                           => n4056);
   U4474 : OAI21_X1 port map( B1 => n5875, B2 => n5888, A => n5744, ZN => n5887
                           );
   U4475 : MUX2_X1 port map( A => REGISTERS_7_63_port, B => n5810, S => n69, Z 
                           => n4055);
   U4476 : MUX2_X1 port map( A => REGISTERS_7_62_port, B => n5812, S => n69, Z 
                           => n4054);
   U4477 : MUX2_X1 port map( A => REGISTERS_7_61_port, B => n5813, S => n69, Z 
                           => n4053);
   U4478 : MUX2_X1 port map( A => REGISTERS_7_60_port, B => n5814, S => n69, Z 
                           => n4052);
   U4479 : MUX2_X1 port map( A => REGISTERS_7_59_port, B => n5815, S => n69, Z 
                           => n4051);
   U4480 : MUX2_X1 port map( A => REGISTERS_7_58_port, B => n5816, S => n69, Z 
                           => n4050);
   U4481 : MUX2_X1 port map( A => REGISTERS_7_57_port, B => n5817, S => n69, Z 
                           => n4049);
   U4482 : MUX2_X1 port map( A => REGISTERS_7_56_port, B => n5818, S => n69, Z 
                           => n4048);
   U4483 : MUX2_X1 port map( A => REGISTERS_7_55_port, B => n5819, S => n69, Z 
                           => n4047);
   U4484 : MUX2_X1 port map( A => REGISTERS_7_54_port, B => n5820, S => n69, Z 
                           => n4046);
   U4485 : MUX2_X1 port map( A => REGISTERS_7_53_port, B => n5821, S => n69, Z 
                           => n4045);
   U4486 : MUX2_X1 port map( A => REGISTERS_7_52_port, B => n5822, S => n69, Z 
                           => n4044);
   U4487 : MUX2_X1 port map( A => REGISTERS_7_51_port, B => n5823, S => n69, Z 
                           => n4043);
   U4488 : MUX2_X1 port map( A => REGISTERS_7_50_port, B => n5824, S => n69, Z 
                           => n4042);
   U4489 : MUX2_X1 port map( A => REGISTERS_7_49_port, B => n5825, S => n69, Z 
                           => n4041);
   U4490 : MUX2_X1 port map( A => REGISTERS_7_48_port, B => n5826, S => n69, Z 
                           => n4040);
   U4491 : MUX2_X1 port map( A => REGISTERS_7_47_port, B => n5827, S => n69, Z 
                           => n4039);
   U4492 : MUX2_X1 port map( A => REGISTERS_7_46_port, B => n5828, S => n69, Z 
                           => n4038);
   U4493 : MUX2_X1 port map( A => REGISTERS_7_45_port, B => n5829, S => n69, Z 
                           => n4037);
   U4494 : MUX2_X1 port map( A => REGISTERS_7_44_port, B => n5830, S => n69, Z 
                           => n4036);
   U4495 : MUX2_X1 port map( A => REGISTERS_7_43_port, B => n5831, S => n69, Z 
                           => n4035);
   U4496 : MUX2_X1 port map( A => REGISTERS_7_42_port, B => n5832, S => n69, Z 
                           => n4034);
   U4497 : MUX2_X1 port map( A => REGISTERS_7_41_port, B => n5833, S => n69, Z 
                           => n4033);
   U4498 : MUX2_X1 port map( A => REGISTERS_7_40_port, B => n5834, S => n69, Z 
                           => n4032);
   U4499 : MUX2_X1 port map( A => REGISTERS_7_39_port, B => n5835, S => n69, Z 
                           => n4031);
   U4500 : MUX2_X1 port map( A => REGISTERS_7_38_port, B => n5836, S => n69, Z 
                           => n4030);
   U4501 : MUX2_X1 port map( A => REGISTERS_7_37_port, B => n5837, S => n69, Z 
                           => n4029);
   U4502 : MUX2_X1 port map( A => REGISTERS_7_36_port, B => n5838, S => n69, Z 
                           => n4028);
   U4503 : MUX2_X1 port map( A => REGISTERS_7_35_port, B => n5839, S => n69, Z 
                           => n4027);
   U4504 : MUX2_X1 port map( A => REGISTERS_7_34_port, B => n5840, S => n69, Z 
                           => n4026);
   U4505 : MUX2_X1 port map( A => REGISTERS_7_33_port, B => n5841, S => n69, Z 
                           => n4025);
   U4506 : MUX2_X1 port map( A => REGISTERS_7_32_port, B => n5842, S => n69, Z 
                           => n4024);
   U4507 : MUX2_X1 port map( A => REGISTERS_7_31_port, B => n5843, S => n69, Z 
                           => n4023);
   U4508 : MUX2_X1 port map( A => REGISTERS_7_30_port, B => n5844, S => n69, Z 
                           => n4022);
   U4509 : MUX2_X1 port map( A => REGISTERS_7_29_port, B => n5845, S => n69, Z 
                           => n4021);
   U4510 : MUX2_X1 port map( A => REGISTERS_7_28_port, B => n5846, S => n69, Z 
                           => n4020);
   U4511 : MUX2_X1 port map( A => REGISTERS_7_27_port, B => n5847, S => n69, Z 
                           => n4019);
   U4512 : MUX2_X1 port map( A => REGISTERS_7_26_port, B => n5848, S => n69, Z 
                           => n4018);
   U4513 : MUX2_X1 port map( A => REGISTERS_7_25_port, B => n5849, S => n69, Z 
                           => n4017);
   U4514 : MUX2_X1 port map( A => REGISTERS_7_24_port, B => n5850, S => n69, Z 
                           => n4016);
   U4515 : MUX2_X1 port map( A => REGISTERS_7_23_port, B => n5851, S => n69, Z 
                           => n4015);
   U4516 : MUX2_X1 port map( A => REGISTERS_7_22_port, B => n5852, S => n69, Z 
                           => n4014);
   U4517 : MUX2_X1 port map( A => REGISTERS_7_21_port, B => n5853, S => n69, Z 
                           => n4013);
   U4518 : MUX2_X1 port map( A => REGISTERS_7_20_port, B => n5854, S => n69, Z 
                           => n4012);
   U4519 : MUX2_X1 port map( A => REGISTERS_7_19_port, B => n5855, S => n69, Z 
                           => n4011);
   U4520 : MUX2_X1 port map( A => REGISTERS_7_18_port, B => n5856, S => n69, Z 
                           => n4010);
   U4521 : MUX2_X1 port map( A => REGISTERS_7_17_port, B => n5857, S => n69, Z 
                           => n4009);
   U4522 : MUX2_X1 port map( A => REGISTERS_7_16_port, B => n5858, S => n69, Z 
                           => n4008);
   U4523 : MUX2_X1 port map( A => REGISTERS_7_15_port, B => n5859, S => n69, Z 
                           => n4007);
   U4524 : MUX2_X1 port map( A => REGISTERS_7_14_port, B => n5860, S => n69, Z 
                           => n4006);
   U4525 : MUX2_X1 port map( A => REGISTERS_7_13_port, B => n5861, S => n69, Z 
                           => n4005);
   U4526 : MUX2_X1 port map( A => REGISTERS_7_12_port, B => n5862, S => n69, Z 
                           => n4004);
   U4527 : MUX2_X1 port map( A => REGISTERS_7_11_port, B => n5863, S => n69, Z 
                           => n4003);
   U4528 : MUX2_X1 port map( A => REGISTERS_7_10_port, B => n5864, S => n69, Z 
                           => n4002);
   U4529 : MUX2_X1 port map( A => REGISTERS_7_9_port, B => n5865, S => n69, Z 
                           => n4001);
   U4530 : MUX2_X1 port map( A => REGISTERS_7_8_port, B => n5866, S => n69, Z 
                           => n4000);
   U4531 : MUX2_X1 port map( A => REGISTERS_7_7_port, B => n5867, S => n69, Z 
                           => n3999);
   U4532 : MUX2_X1 port map( A => REGISTERS_7_6_port, B => n5868, S => n69, Z 
                           => n3998);
   U4533 : MUX2_X1 port map( A => REGISTERS_7_5_port, B => n5869, S => n69, Z 
                           => n3997);
   U4534 : MUX2_X1 port map( A => REGISTERS_7_4_port, B => n5870, S => n69, Z 
                           => n3996);
   U4535 : MUX2_X1 port map( A => REGISTERS_7_3_port, B => n5871, S => n69, Z 
                           => n3995);
   U4536 : MUX2_X1 port map( A => REGISTERS_7_2_port, B => n5872, S => n69, Z 
                           => n3994);
   U4537 : MUX2_X1 port map( A => REGISTERS_7_1_port, B => n5873, S => n69, Z 
                           => n3993);
   U4538 : MUX2_X1 port map( A => REGISTERS_7_0_port, B => n5874, S => n69, Z 
                           => n3992);
   U4539 : OAI21_X1 port map( B1 => n5875, B2 => n5890, A => n5744, ZN => n5889
                           );
   U4540 : NAND3_X1 port map( A1 => n5891, A2 => n5892, A3 => n5893, ZN => 
                           n5875);
   U4541 : MUX2_X1 port map( A => REGISTERS_8_63_port, B => n5810, S => n71, Z 
                           => n3991);
   U4542 : MUX2_X1 port map( A => REGISTERS_8_62_port, B => n5812, S => n71, Z 
                           => n3990);
   U4543 : MUX2_X1 port map( A => REGISTERS_8_61_port, B => n5813, S => n71, Z 
                           => n3989);
   U4544 : MUX2_X1 port map( A => REGISTERS_8_60_port, B => n5814, S => n71, Z 
                           => n3988);
   U4545 : MUX2_X1 port map( A => REGISTERS_8_59_port, B => n5815, S => n71, Z 
                           => n3987);
   U4546 : MUX2_X1 port map( A => REGISTERS_8_58_port, B => n5816, S => n71, Z 
                           => n3986);
   U4547 : MUX2_X1 port map( A => REGISTERS_8_57_port, B => n5817, S => n71, Z 
                           => n3985);
   U4548 : MUX2_X1 port map( A => REGISTERS_8_56_port, B => n5818, S => n71, Z 
                           => n3984);
   U4549 : MUX2_X1 port map( A => REGISTERS_8_55_port, B => n5819, S => n71, Z 
                           => n3983);
   U4550 : MUX2_X1 port map( A => REGISTERS_8_54_port, B => n5820, S => n71, Z 
                           => n3982);
   U4551 : MUX2_X1 port map( A => REGISTERS_8_53_port, B => n5821, S => n71, Z 
                           => n3981);
   U4552 : MUX2_X1 port map( A => REGISTERS_8_52_port, B => n5822, S => n71, Z 
                           => n3980);
   U4553 : MUX2_X1 port map( A => REGISTERS_8_51_port, B => n5823, S => n71, Z 
                           => n3979);
   U4554 : MUX2_X1 port map( A => REGISTERS_8_50_port, B => n5824, S => n71, Z 
                           => n3978);
   U4555 : MUX2_X1 port map( A => REGISTERS_8_49_port, B => n5825, S => n71, Z 
                           => n3977);
   U4556 : MUX2_X1 port map( A => REGISTERS_8_48_port, B => n5826, S => n71, Z 
                           => n3976);
   U4557 : MUX2_X1 port map( A => REGISTERS_8_47_port, B => n5827, S => n71, Z 
                           => n3975);
   U4558 : MUX2_X1 port map( A => REGISTERS_8_46_port, B => n5828, S => n71, Z 
                           => n3974);
   U4559 : MUX2_X1 port map( A => REGISTERS_8_45_port, B => n5829, S => n71, Z 
                           => n3973);
   U4560 : MUX2_X1 port map( A => REGISTERS_8_44_port, B => n5830, S => n71, Z 
                           => n3972);
   U4561 : MUX2_X1 port map( A => REGISTERS_8_43_port, B => n5831, S => n71, Z 
                           => n3971);
   U4562 : MUX2_X1 port map( A => REGISTERS_8_42_port, B => n5832, S => n71, Z 
                           => n3970);
   U4563 : MUX2_X1 port map( A => REGISTERS_8_41_port, B => n5833, S => n71, Z 
                           => n3969);
   U4564 : MUX2_X1 port map( A => REGISTERS_8_40_port, B => n5834, S => n71, Z 
                           => n3968);
   U4565 : MUX2_X1 port map( A => REGISTERS_8_39_port, B => n5835, S => n71, Z 
                           => n3967);
   U4566 : MUX2_X1 port map( A => REGISTERS_8_38_port, B => n5836, S => n71, Z 
                           => n3966);
   U4567 : MUX2_X1 port map( A => REGISTERS_8_37_port, B => n5837, S => n71, Z 
                           => n3965);
   U4568 : MUX2_X1 port map( A => REGISTERS_8_36_port, B => n5838, S => n71, Z 
                           => n3964);
   U4569 : MUX2_X1 port map( A => REGISTERS_8_35_port, B => n5839, S => n71, Z 
                           => n3963);
   U4570 : MUX2_X1 port map( A => REGISTERS_8_34_port, B => n5840, S => n71, Z 
                           => n3962);
   U4571 : MUX2_X1 port map( A => REGISTERS_8_33_port, B => n5841, S => n71, Z 
                           => n3961);
   U4572 : MUX2_X1 port map( A => REGISTERS_8_32_port, B => n5842, S => n71, Z 
                           => n3960);
   U4573 : MUX2_X1 port map( A => REGISTERS_8_31_port, B => n5843, S => n71, Z 
                           => n3959);
   U4574 : MUX2_X1 port map( A => REGISTERS_8_30_port, B => n5844, S => n71, Z 
                           => n3958);
   U4575 : MUX2_X1 port map( A => REGISTERS_8_29_port, B => n5845, S => n71, Z 
                           => n3957);
   U4576 : MUX2_X1 port map( A => REGISTERS_8_28_port, B => n5846, S => n71, Z 
                           => n3956);
   U4577 : MUX2_X1 port map( A => REGISTERS_8_27_port, B => n5847, S => n71, Z 
                           => n3955);
   U4578 : MUX2_X1 port map( A => REGISTERS_8_26_port, B => n5848, S => n71, Z 
                           => n3954);
   U4579 : MUX2_X1 port map( A => REGISTERS_8_25_port, B => n5849, S => n71, Z 
                           => n3953);
   U4580 : MUX2_X1 port map( A => REGISTERS_8_24_port, B => n5850, S => n71, Z 
                           => n3952);
   U4581 : MUX2_X1 port map( A => REGISTERS_8_23_port, B => n5851, S => n71, Z 
                           => n3951);
   U4582 : MUX2_X1 port map( A => REGISTERS_8_22_port, B => n5852, S => n71, Z 
                           => n3950);
   U4583 : MUX2_X1 port map( A => REGISTERS_8_21_port, B => n5853, S => n71, Z 
                           => n3949);
   U4584 : MUX2_X1 port map( A => REGISTERS_8_20_port, B => n5854, S => n71, Z 
                           => n3948);
   U4585 : MUX2_X1 port map( A => REGISTERS_8_19_port, B => n5855, S => n71, Z 
                           => n3947);
   U4586 : MUX2_X1 port map( A => REGISTERS_8_18_port, B => n5856, S => n71, Z 
                           => n3946);
   U4587 : MUX2_X1 port map( A => REGISTERS_8_17_port, B => n5857, S => n71, Z 
                           => n3945);
   U4588 : MUX2_X1 port map( A => REGISTERS_8_16_port, B => n5858, S => n71, Z 
                           => n3944);
   U4589 : MUX2_X1 port map( A => REGISTERS_8_15_port, B => n5859, S => n71, Z 
                           => n3943);
   U4590 : MUX2_X1 port map( A => REGISTERS_8_14_port, B => n5860, S => n71, Z 
                           => n3942);
   U4591 : MUX2_X1 port map( A => REGISTERS_8_13_port, B => n5861, S => n71, Z 
                           => n3941);
   U4592 : MUX2_X1 port map( A => REGISTERS_8_12_port, B => n5862, S => n71, Z 
                           => n3940);
   U4593 : MUX2_X1 port map( A => REGISTERS_8_11_port, B => n5863, S => n71, Z 
                           => n3939);
   U4594 : MUX2_X1 port map( A => REGISTERS_8_10_port, B => n5864, S => n71, Z 
                           => n3938);
   U4595 : MUX2_X1 port map( A => REGISTERS_8_9_port, B => n5865, S => n71, Z 
                           => n3937);
   U4596 : MUX2_X1 port map( A => REGISTERS_8_8_port, B => n5866, S => n71, Z 
                           => n3936);
   U4597 : MUX2_X1 port map( A => REGISTERS_8_7_port, B => n5867, S => n71, Z 
                           => n3935);
   U4598 : MUX2_X1 port map( A => REGISTERS_8_6_port, B => n5868, S => n71, Z 
                           => n3934);
   U4599 : MUX2_X1 port map( A => REGISTERS_8_5_port, B => n5869, S => n71, Z 
                           => n3933);
   U4600 : MUX2_X1 port map( A => REGISTERS_8_4_port, B => n5870, S => n71, Z 
                           => n3932);
   U4601 : MUX2_X1 port map( A => REGISTERS_8_3_port, B => n5871, S => n71, Z 
                           => n3931);
   U4602 : MUX2_X1 port map( A => REGISTERS_8_2_port, B => n5872, S => n71, Z 
                           => n3930);
   U4603 : MUX2_X1 port map( A => REGISTERS_8_1_port, B => n5873, S => n71, Z 
                           => n3929);
   U4604 : MUX2_X1 port map( A => REGISTERS_8_0_port, B => n5874, S => n71, Z 
                           => n3928);
   U4605 : OAI21_X1 port map( B1 => n5876, B2 => n5895, A => n5744, ZN => n5894
                           );
   U4606 : MUX2_X1 port map( A => REGISTERS_9_63_port, B => n5810, S => n73, Z 
                           => n3927);
   U4607 : MUX2_X1 port map( A => REGISTERS_9_62_port, B => n5812, S => n73, Z 
                           => n3926);
   U4608 : MUX2_X1 port map( A => REGISTERS_9_61_port, B => n5813, S => n73, Z 
                           => n3925);
   U4609 : MUX2_X1 port map( A => REGISTERS_9_60_port, B => n5814, S => n73, Z 
                           => n3924);
   U4610 : MUX2_X1 port map( A => REGISTERS_9_59_port, B => n5815, S => n73, Z 
                           => n3923);
   U4611 : MUX2_X1 port map( A => REGISTERS_9_58_port, B => n5816, S => n73, Z 
                           => n3922);
   U4612 : MUX2_X1 port map( A => REGISTERS_9_57_port, B => n5817, S => n73, Z 
                           => n3921);
   U4613 : MUX2_X1 port map( A => REGISTERS_9_56_port, B => n5818, S => n73, Z 
                           => n3920);
   U4614 : MUX2_X1 port map( A => REGISTERS_9_55_port, B => n5819, S => n73, Z 
                           => n3919);
   U4615 : MUX2_X1 port map( A => REGISTERS_9_54_port, B => n5820, S => n73, Z 
                           => n3918);
   U4616 : MUX2_X1 port map( A => REGISTERS_9_53_port, B => n5821, S => n73, Z 
                           => n3917);
   U4617 : MUX2_X1 port map( A => REGISTERS_9_52_port, B => n5822, S => n73, Z 
                           => n3916);
   U4618 : MUX2_X1 port map( A => REGISTERS_9_51_port, B => n5823, S => n73, Z 
                           => n3915);
   U4619 : MUX2_X1 port map( A => REGISTERS_9_50_port, B => n5824, S => n73, Z 
                           => n3914);
   U4620 : MUX2_X1 port map( A => REGISTERS_9_49_port, B => n5825, S => n73, Z 
                           => n3913);
   U4621 : MUX2_X1 port map( A => REGISTERS_9_48_port, B => n5826, S => n73, Z 
                           => n3912);
   U4622 : MUX2_X1 port map( A => REGISTERS_9_47_port, B => n5827, S => n73, Z 
                           => n3911);
   U4623 : MUX2_X1 port map( A => REGISTERS_9_46_port, B => n5828, S => n73, Z 
                           => n3910);
   U4624 : MUX2_X1 port map( A => REGISTERS_9_45_port, B => n5829, S => n73, Z 
                           => n3909);
   U4625 : MUX2_X1 port map( A => REGISTERS_9_44_port, B => n5830, S => n73, Z 
                           => n3908);
   U4626 : MUX2_X1 port map( A => REGISTERS_9_43_port, B => n5831, S => n73, Z 
                           => n3907);
   U4627 : MUX2_X1 port map( A => REGISTERS_9_42_port, B => n5832, S => n73, Z 
                           => n3906);
   U4628 : MUX2_X1 port map( A => REGISTERS_9_41_port, B => n5833, S => n73, Z 
                           => n3905);
   U4629 : MUX2_X1 port map( A => REGISTERS_9_40_port, B => n5834, S => n73, Z 
                           => n3904);
   U4630 : MUX2_X1 port map( A => REGISTERS_9_39_port, B => n5835, S => n73, Z 
                           => n3903);
   U4631 : MUX2_X1 port map( A => REGISTERS_9_38_port, B => n5836, S => n73, Z 
                           => n3902);
   U4632 : MUX2_X1 port map( A => REGISTERS_9_37_port, B => n5837, S => n73, Z 
                           => n3901);
   U4633 : MUX2_X1 port map( A => REGISTERS_9_36_port, B => n5838, S => n73, Z 
                           => n3900);
   U4634 : MUX2_X1 port map( A => REGISTERS_9_35_port, B => n5839, S => n73, Z 
                           => n3899);
   U4635 : MUX2_X1 port map( A => REGISTERS_9_34_port, B => n5840, S => n73, Z 
                           => n3898);
   U4636 : MUX2_X1 port map( A => REGISTERS_9_33_port, B => n5841, S => n73, Z 
                           => n3897);
   U4637 : MUX2_X1 port map( A => REGISTERS_9_32_port, B => n5842, S => n73, Z 
                           => n3896);
   U4638 : MUX2_X1 port map( A => REGISTERS_9_31_port, B => n5843, S => n73, Z 
                           => n3895);
   U4639 : MUX2_X1 port map( A => REGISTERS_9_30_port, B => n5844, S => n73, Z 
                           => n3894);
   U4640 : MUX2_X1 port map( A => REGISTERS_9_29_port, B => n5845, S => n73, Z 
                           => n3893);
   U4641 : MUX2_X1 port map( A => REGISTERS_9_28_port, B => n5846, S => n73, Z 
                           => n3892);
   U4642 : MUX2_X1 port map( A => REGISTERS_9_27_port, B => n5847, S => n73, Z 
                           => n3891);
   U4643 : MUX2_X1 port map( A => REGISTERS_9_26_port, B => n5848, S => n73, Z 
                           => n3890);
   U4644 : MUX2_X1 port map( A => REGISTERS_9_25_port, B => n5849, S => n73, Z 
                           => n3889);
   U4645 : MUX2_X1 port map( A => REGISTERS_9_24_port, B => n5850, S => n73, Z 
                           => n3888);
   U4646 : MUX2_X1 port map( A => REGISTERS_9_23_port, B => n5851, S => n73, Z 
                           => n3887);
   U4647 : MUX2_X1 port map( A => REGISTERS_9_22_port, B => n5852, S => n73, Z 
                           => n3886);
   U4648 : MUX2_X1 port map( A => REGISTERS_9_21_port, B => n5853, S => n73, Z 
                           => n3885);
   U4649 : MUX2_X1 port map( A => REGISTERS_9_20_port, B => n5854, S => n73, Z 
                           => n3884);
   U4650 : MUX2_X1 port map( A => REGISTERS_9_19_port, B => n5855, S => n73, Z 
                           => n3883);
   U4651 : MUX2_X1 port map( A => REGISTERS_9_18_port, B => n5856, S => n73, Z 
                           => n3882);
   U4652 : MUX2_X1 port map( A => REGISTERS_9_17_port, B => n5857, S => n73, Z 
                           => n3881);
   U4653 : MUX2_X1 port map( A => REGISTERS_9_16_port, B => n5858, S => n73, Z 
                           => n3880);
   U4654 : MUX2_X1 port map( A => REGISTERS_9_15_port, B => n5859, S => n73, Z 
                           => n3879);
   U4655 : MUX2_X1 port map( A => REGISTERS_9_14_port, B => n5860, S => n73, Z 
                           => n3878);
   U4656 : MUX2_X1 port map( A => REGISTERS_9_13_port, B => n5861, S => n73, Z 
                           => n3877);
   U4657 : MUX2_X1 port map( A => REGISTERS_9_12_port, B => n5862, S => n73, Z 
                           => n3876);
   U4658 : MUX2_X1 port map( A => REGISTERS_9_11_port, B => n5863, S => n73, Z 
                           => n3875);
   U4659 : MUX2_X1 port map( A => REGISTERS_9_10_port, B => n5864, S => n73, Z 
                           => n3874);
   U4660 : MUX2_X1 port map( A => REGISTERS_9_9_port, B => n5865, S => n73, Z 
                           => n3873);
   U4661 : MUX2_X1 port map( A => REGISTERS_9_8_port, B => n5866, S => n73, Z 
                           => n3872);
   U4662 : MUX2_X1 port map( A => REGISTERS_9_7_port, B => n5867, S => n73, Z 
                           => n3871);
   U4663 : MUX2_X1 port map( A => REGISTERS_9_6_port, B => n5868, S => n73, Z 
                           => n3870);
   U4664 : MUX2_X1 port map( A => REGISTERS_9_5_port, B => n5869, S => n73, Z 
                           => n3869);
   U4665 : MUX2_X1 port map( A => REGISTERS_9_4_port, B => n5870, S => n73, Z 
                           => n3868);
   U4666 : MUX2_X1 port map( A => REGISTERS_9_3_port, B => n5871, S => n73, Z 
                           => n3867);
   U4667 : MUX2_X1 port map( A => REGISTERS_9_2_port, B => n5872, S => n73, Z 
                           => n3866);
   U4668 : MUX2_X1 port map( A => REGISTERS_9_1_port, B => n5873, S => n73, Z 
                           => n3865);
   U4669 : MUX2_X1 port map( A => REGISTERS_9_0_port, B => n5874, S => n73, Z 
                           => n3864);
   U4670 : OAI21_X1 port map( B1 => n5878, B2 => n5895, A => n5744, ZN => n5896
                           );
   U4671 : MUX2_X1 port map( A => REGISTERS_10_63_port, B => n5810, S => n75, Z
                           => n3863);
   U4672 : MUX2_X1 port map( A => REGISTERS_10_62_port, B => n5812, S => n75, Z
                           => n3862);
   U4673 : MUX2_X1 port map( A => REGISTERS_10_61_port, B => n5813, S => n75, Z
                           => n3861);
   U4674 : MUX2_X1 port map( A => REGISTERS_10_60_port, B => n5814, S => n75, Z
                           => n3860);
   U4675 : MUX2_X1 port map( A => REGISTERS_10_59_port, B => n5815, S => n75, Z
                           => n3859);
   U4676 : MUX2_X1 port map( A => REGISTERS_10_58_port, B => n5816, S => n75, Z
                           => n3858);
   U4677 : MUX2_X1 port map( A => REGISTERS_10_57_port, B => n5817, S => n75, Z
                           => n3857);
   U4678 : MUX2_X1 port map( A => REGISTERS_10_56_port, B => n5818, S => n75, Z
                           => n3856);
   U4679 : MUX2_X1 port map( A => REGISTERS_10_55_port, B => n5819, S => n75, Z
                           => n3855);
   U4680 : MUX2_X1 port map( A => REGISTERS_10_54_port, B => n5820, S => n75, Z
                           => n3854);
   U4681 : MUX2_X1 port map( A => REGISTERS_10_53_port, B => n5821, S => n75, Z
                           => n3853);
   U4682 : MUX2_X1 port map( A => REGISTERS_10_52_port, B => n5822, S => n75, Z
                           => n3852);
   U4683 : MUX2_X1 port map( A => REGISTERS_10_51_port, B => n5823, S => n75, Z
                           => n3851);
   U4684 : MUX2_X1 port map( A => REGISTERS_10_50_port, B => n5824, S => n75, Z
                           => n3850);
   U4685 : MUX2_X1 port map( A => REGISTERS_10_49_port, B => n5825, S => n75, Z
                           => n3849);
   U4686 : MUX2_X1 port map( A => REGISTERS_10_48_port, B => n5826, S => n75, Z
                           => n3848);
   U4687 : MUX2_X1 port map( A => REGISTERS_10_47_port, B => n5827, S => n75, Z
                           => n3847);
   U4688 : MUX2_X1 port map( A => REGISTERS_10_46_port, B => n5828, S => n75, Z
                           => n3846);
   U4689 : MUX2_X1 port map( A => REGISTERS_10_45_port, B => n5829, S => n75, Z
                           => n3845);
   U4690 : MUX2_X1 port map( A => REGISTERS_10_44_port, B => n5830, S => n75, Z
                           => n3844);
   U4691 : MUX2_X1 port map( A => REGISTERS_10_43_port, B => n5831, S => n75, Z
                           => n3843);
   U4692 : MUX2_X1 port map( A => REGISTERS_10_42_port, B => n5832, S => n75, Z
                           => n3842);
   U4693 : MUX2_X1 port map( A => REGISTERS_10_41_port, B => n5833, S => n75, Z
                           => n3841);
   U4694 : MUX2_X1 port map( A => REGISTERS_10_40_port, B => n5834, S => n75, Z
                           => n3840);
   U4695 : MUX2_X1 port map( A => REGISTERS_10_39_port, B => n5835, S => n75, Z
                           => n3839);
   U4696 : MUX2_X1 port map( A => REGISTERS_10_38_port, B => n5836, S => n75, Z
                           => n3838);
   U4697 : MUX2_X1 port map( A => REGISTERS_10_37_port, B => n5837, S => n75, Z
                           => n3837);
   U4698 : MUX2_X1 port map( A => REGISTERS_10_36_port, B => n5838, S => n75, Z
                           => n3836);
   U4699 : MUX2_X1 port map( A => REGISTERS_10_35_port, B => n5839, S => n75, Z
                           => n3835);
   U4700 : MUX2_X1 port map( A => REGISTERS_10_34_port, B => n5840, S => n75, Z
                           => n3834);
   U4701 : MUX2_X1 port map( A => REGISTERS_10_33_port, B => n5841, S => n75, Z
                           => n3833);
   U4702 : MUX2_X1 port map( A => REGISTERS_10_32_port, B => n5842, S => n75, Z
                           => n3832);
   U4703 : MUX2_X1 port map( A => REGISTERS_10_31_port, B => n5843, S => n75, Z
                           => n3831);
   U4704 : MUX2_X1 port map( A => REGISTERS_10_30_port, B => n5844, S => n75, Z
                           => n3830);
   U4705 : MUX2_X1 port map( A => REGISTERS_10_29_port, B => n5845, S => n75, Z
                           => n3829);
   U4706 : MUX2_X1 port map( A => REGISTERS_10_28_port, B => n5846, S => n75, Z
                           => n3828);
   U4707 : MUX2_X1 port map( A => REGISTERS_10_27_port, B => n5847, S => n75, Z
                           => n3827);
   U4708 : MUX2_X1 port map( A => REGISTERS_10_26_port, B => n5848, S => n75, Z
                           => n3826);
   U4709 : MUX2_X1 port map( A => REGISTERS_10_25_port, B => n5849, S => n75, Z
                           => n3825);
   U4710 : MUX2_X1 port map( A => REGISTERS_10_24_port, B => n5850, S => n75, Z
                           => n3824);
   U4711 : MUX2_X1 port map( A => REGISTERS_10_23_port, B => n5851, S => n75, Z
                           => n3823);
   U4712 : MUX2_X1 port map( A => REGISTERS_10_22_port, B => n5852, S => n75, Z
                           => n3822);
   U4713 : MUX2_X1 port map( A => REGISTERS_10_21_port, B => n5853, S => n75, Z
                           => n3821);
   U4714 : MUX2_X1 port map( A => REGISTERS_10_20_port, B => n5854, S => n75, Z
                           => n3820);
   U4715 : MUX2_X1 port map( A => REGISTERS_10_19_port, B => n5855, S => n75, Z
                           => n3819);
   U4716 : MUX2_X1 port map( A => REGISTERS_10_18_port, B => n5856, S => n75, Z
                           => n3818);
   U4717 : MUX2_X1 port map( A => REGISTERS_10_17_port, B => n5857, S => n75, Z
                           => n3817);
   U4718 : MUX2_X1 port map( A => REGISTERS_10_16_port, B => n5858, S => n75, Z
                           => n3816);
   U4719 : MUX2_X1 port map( A => REGISTERS_10_15_port, B => n5859, S => n75, Z
                           => n3815);
   U4720 : MUX2_X1 port map( A => REGISTERS_10_14_port, B => n5860, S => n75, Z
                           => n3814);
   U4721 : MUX2_X1 port map( A => REGISTERS_10_13_port, B => n5861, S => n75, Z
                           => n3813);
   U4722 : MUX2_X1 port map( A => REGISTERS_10_12_port, B => n5862, S => n75, Z
                           => n3812);
   U4723 : MUX2_X1 port map( A => REGISTERS_10_11_port, B => n5863, S => n75, Z
                           => n3811);
   U4724 : MUX2_X1 port map( A => REGISTERS_10_10_port, B => n5864, S => n75, Z
                           => n3810);
   U4725 : MUX2_X1 port map( A => REGISTERS_10_9_port, B => n5865, S => n75, Z 
                           => n3809);
   U4726 : MUX2_X1 port map( A => REGISTERS_10_8_port, B => n5866, S => n75, Z 
                           => n3808);
   U4727 : MUX2_X1 port map( A => REGISTERS_10_7_port, B => n5867, S => n75, Z 
                           => n3807);
   U4728 : MUX2_X1 port map( A => REGISTERS_10_6_port, B => n5868, S => n75, Z 
                           => n3806);
   U4729 : MUX2_X1 port map( A => REGISTERS_10_5_port, B => n5869, S => n75, Z 
                           => n3805);
   U4730 : MUX2_X1 port map( A => REGISTERS_10_4_port, B => n5870, S => n75, Z 
                           => n3804);
   U4731 : MUX2_X1 port map( A => REGISTERS_10_3_port, B => n5871, S => n75, Z 
                           => n3803);
   U4732 : MUX2_X1 port map( A => REGISTERS_10_2_port, B => n5872, S => n75, Z 
                           => n3802);
   U4733 : MUX2_X1 port map( A => REGISTERS_10_1_port, B => n5873, S => n75, Z 
                           => n3801);
   U4734 : MUX2_X1 port map( A => REGISTERS_10_0_port, B => n5874, S => n75, Z 
                           => n3800);
   U4735 : OAI21_X1 port map( B1 => n5880, B2 => n5895, A => n5744, ZN => n5897
                           );
   U4736 : MUX2_X1 port map( A => REGISTERS_11_63_port, B => n5810, S => n61, Z
                           => n3799);
   U4737 : MUX2_X1 port map( A => REGISTERS_11_62_port, B => n5812, S => n61, Z
                           => n3798);
   U4738 : MUX2_X1 port map( A => REGISTERS_11_61_port, B => n5813, S => n61, Z
                           => n3797);
   U4739 : MUX2_X1 port map( A => REGISTERS_11_60_port, B => n5814, S => n61, Z
                           => n3796);
   U4740 : MUX2_X1 port map( A => REGISTERS_11_59_port, B => n5815, S => n61, Z
                           => n3795);
   U4741 : MUX2_X1 port map( A => REGISTERS_11_58_port, B => n5816, S => n61, Z
                           => n3794);
   U4742 : MUX2_X1 port map( A => REGISTERS_11_57_port, B => n5817, S => n61, Z
                           => n3793);
   U4743 : MUX2_X1 port map( A => REGISTERS_11_56_port, B => n5818, S => n61, Z
                           => n3792);
   U4744 : MUX2_X1 port map( A => REGISTERS_11_55_port, B => n5819, S => n61, Z
                           => n3791);
   U4745 : MUX2_X1 port map( A => REGISTERS_11_54_port, B => n5820, S => n61, Z
                           => n3790);
   U4746 : MUX2_X1 port map( A => REGISTERS_11_53_port, B => n5821, S => n61, Z
                           => n3789);
   U4747 : MUX2_X1 port map( A => REGISTERS_11_52_port, B => n5822, S => n61, Z
                           => n3788);
   U4748 : MUX2_X1 port map( A => REGISTERS_11_51_port, B => n5823, S => n61, Z
                           => n3787);
   U4749 : MUX2_X1 port map( A => REGISTERS_11_50_port, B => n5824, S => n61, Z
                           => n3786);
   U4750 : MUX2_X1 port map( A => REGISTERS_11_49_port, B => n5825, S => n61, Z
                           => n3785);
   U4751 : MUX2_X1 port map( A => REGISTERS_11_48_port, B => n5826, S => n61, Z
                           => n3784);
   U4752 : MUX2_X1 port map( A => REGISTERS_11_47_port, B => n5827, S => n61, Z
                           => n3783);
   U4753 : MUX2_X1 port map( A => REGISTERS_11_46_port, B => n5828, S => n61, Z
                           => n3782);
   U4754 : MUX2_X1 port map( A => REGISTERS_11_45_port, B => n5829, S => n61, Z
                           => n3781);
   U4755 : MUX2_X1 port map( A => REGISTERS_11_44_port, B => n5830, S => n61, Z
                           => n3780);
   U4756 : MUX2_X1 port map( A => REGISTERS_11_43_port, B => n5831, S => n61, Z
                           => n3779);
   U4757 : MUX2_X1 port map( A => REGISTERS_11_42_port, B => n5832, S => n61, Z
                           => n3778);
   U4758 : MUX2_X1 port map( A => REGISTERS_11_41_port, B => n5833, S => n61, Z
                           => n3777);
   U4759 : MUX2_X1 port map( A => REGISTERS_11_40_port, B => n5834, S => n61, Z
                           => n3776);
   U4760 : MUX2_X1 port map( A => REGISTERS_11_39_port, B => n5835, S => n61, Z
                           => n3775);
   U4761 : MUX2_X1 port map( A => REGISTERS_11_38_port, B => n5836, S => n61, Z
                           => n3774);
   U4762 : MUX2_X1 port map( A => REGISTERS_11_37_port, B => n5837, S => n61, Z
                           => n3773);
   U4763 : MUX2_X1 port map( A => REGISTERS_11_36_port, B => n5838, S => n61, Z
                           => n3772);
   U4764 : MUX2_X1 port map( A => REGISTERS_11_35_port, B => n5839, S => n61, Z
                           => n3771);
   U4765 : MUX2_X1 port map( A => REGISTERS_11_34_port, B => n5840, S => n61, Z
                           => n3770);
   U4766 : MUX2_X1 port map( A => REGISTERS_11_33_port, B => n5841, S => n61, Z
                           => n3769);
   U4767 : MUX2_X1 port map( A => REGISTERS_11_32_port, B => n5842, S => n61, Z
                           => n3768);
   U4768 : MUX2_X1 port map( A => REGISTERS_11_31_port, B => n5843, S => n61, Z
                           => n3767);
   U4769 : MUX2_X1 port map( A => REGISTERS_11_30_port, B => n5844, S => n61, Z
                           => n3766);
   U4770 : MUX2_X1 port map( A => REGISTERS_11_29_port, B => n5845, S => n61, Z
                           => n3765);
   U4771 : MUX2_X1 port map( A => REGISTERS_11_28_port, B => n5846, S => n61, Z
                           => n3764);
   U4772 : MUX2_X1 port map( A => REGISTERS_11_27_port, B => n5847, S => n61, Z
                           => n3763);
   U4773 : MUX2_X1 port map( A => REGISTERS_11_26_port, B => n5848, S => n61, Z
                           => n3762);
   U4774 : MUX2_X1 port map( A => REGISTERS_11_25_port, B => n5849, S => n61, Z
                           => n3761);
   U4775 : MUX2_X1 port map( A => REGISTERS_11_24_port, B => n5850, S => n61, Z
                           => n3760);
   U4776 : MUX2_X1 port map( A => REGISTERS_11_23_port, B => n5851, S => n61, Z
                           => n3759);
   U4777 : MUX2_X1 port map( A => REGISTERS_11_22_port, B => n5852, S => n61, Z
                           => n3758);
   U4778 : MUX2_X1 port map( A => REGISTERS_11_21_port, B => n5853, S => n61, Z
                           => n3757);
   U4779 : MUX2_X1 port map( A => REGISTERS_11_20_port, B => n5854, S => n61, Z
                           => n3756);
   U4780 : MUX2_X1 port map( A => REGISTERS_11_19_port, B => n5855, S => n61, Z
                           => n3755);
   U4781 : MUX2_X1 port map( A => REGISTERS_11_18_port, B => n5856, S => n61, Z
                           => n3754);
   U4782 : MUX2_X1 port map( A => REGISTERS_11_17_port, B => n5857, S => n61, Z
                           => n3753);
   U4783 : MUX2_X1 port map( A => REGISTERS_11_16_port, B => n5858, S => n61, Z
                           => n3752);
   U4784 : MUX2_X1 port map( A => REGISTERS_11_15_port, B => n5859, S => n61, Z
                           => n3751);
   U4785 : MUX2_X1 port map( A => REGISTERS_11_14_port, B => n5860, S => n61, Z
                           => n3750);
   U4786 : MUX2_X1 port map( A => REGISTERS_11_13_port, B => n5861, S => n61, Z
                           => n3749);
   U4787 : MUX2_X1 port map( A => REGISTERS_11_12_port, B => n5862, S => n61, Z
                           => n3748);
   U4788 : MUX2_X1 port map( A => REGISTERS_11_11_port, B => n5863, S => n61, Z
                           => n3747);
   U4789 : MUX2_X1 port map( A => REGISTERS_11_10_port, B => n5864, S => n61, Z
                           => n3746);
   U4790 : MUX2_X1 port map( A => REGISTERS_11_9_port, B => n5865, S => n61, Z 
                           => n3745);
   U4791 : MUX2_X1 port map( A => REGISTERS_11_8_port, B => n5866, S => n61, Z 
                           => n3744);
   U4792 : MUX2_X1 port map( A => REGISTERS_11_7_port, B => n5867, S => n61, Z 
                           => n3743);
   U4793 : MUX2_X1 port map( A => REGISTERS_11_6_port, B => n5868, S => n61, Z 
                           => n3742);
   U4794 : MUX2_X1 port map( A => REGISTERS_11_5_port, B => n5869, S => n61, Z 
                           => n3741);
   U4795 : MUX2_X1 port map( A => REGISTERS_11_4_port, B => n5870, S => n61, Z 
                           => n3740);
   U4796 : MUX2_X1 port map( A => REGISTERS_11_3_port, B => n5871, S => n61, Z 
                           => n3739);
   U4797 : MUX2_X1 port map( A => REGISTERS_11_2_port, B => n5872, S => n61, Z 
                           => n3738);
   U4798 : MUX2_X1 port map( A => REGISTERS_11_1_port, B => n5873, S => n61, Z 
                           => n3737);
   U4799 : MUX2_X1 port map( A => REGISTERS_11_0_port, B => n5874, S => n61, Z 
                           => n3736);
   U4800 : OAI21_X1 port map( B1 => n5882, B2 => n5895, A => n5744, ZN => n5898
                           );
   U4801 : MUX2_X1 port map( A => REGISTERS_12_63_port, B => n5810, S => n63, Z
                           => n3735);
   U4802 : MUX2_X1 port map( A => REGISTERS_12_62_port, B => n5812, S => n63, Z
                           => n3734);
   U4803 : MUX2_X1 port map( A => REGISTERS_12_61_port, B => n5813, S => n63, Z
                           => n3733);
   U4804 : MUX2_X1 port map( A => REGISTERS_12_60_port, B => n5814, S => n63, Z
                           => n3732);
   U4805 : MUX2_X1 port map( A => REGISTERS_12_59_port, B => n5815, S => n63, Z
                           => n3731);
   U4806 : MUX2_X1 port map( A => REGISTERS_12_58_port, B => n5816, S => n63, Z
                           => n3730);
   U4807 : MUX2_X1 port map( A => REGISTERS_12_57_port, B => n5817, S => n63, Z
                           => n3729);
   U4808 : MUX2_X1 port map( A => REGISTERS_12_56_port, B => n5818, S => n63, Z
                           => n3728);
   U4809 : MUX2_X1 port map( A => REGISTERS_12_55_port, B => n5819, S => n63, Z
                           => n3727);
   U4810 : MUX2_X1 port map( A => REGISTERS_12_54_port, B => n5820, S => n63, Z
                           => n3726);
   U4811 : MUX2_X1 port map( A => REGISTERS_12_53_port, B => n5821, S => n63, Z
                           => n3725);
   U4812 : MUX2_X1 port map( A => REGISTERS_12_52_port, B => n5822, S => n63, Z
                           => n3724);
   U4813 : MUX2_X1 port map( A => REGISTERS_12_51_port, B => n5823, S => n63, Z
                           => n3723);
   U4814 : MUX2_X1 port map( A => REGISTERS_12_50_port, B => n5824, S => n63, Z
                           => n3722);
   U4815 : MUX2_X1 port map( A => REGISTERS_12_49_port, B => n5825, S => n63, Z
                           => n3721);
   U4816 : MUX2_X1 port map( A => REGISTERS_12_48_port, B => n5826, S => n63, Z
                           => n3720);
   U4817 : MUX2_X1 port map( A => REGISTERS_12_47_port, B => n5827, S => n63, Z
                           => n3719);
   U4818 : MUX2_X1 port map( A => REGISTERS_12_46_port, B => n5828, S => n63, Z
                           => n3718);
   U4819 : MUX2_X1 port map( A => REGISTERS_12_45_port, B => n5829, S => n63, Z
                           => n3717);
   U4820 : MUX2_X1 port map( A => REGISTERS_12_44_port, B => n5830, S => n63, Z
                           => n3716);
   U4821 : MUX2_X1 port map( A => REGISTERS_12_43_port, B => n5831, S => n63, Z
                           => n3715);
   U4822 : MUX2_X1 port map( A => REGISTERS_12_42_port, B => n5832, S => n63, Z
                           => n3714);
   U4823 : MUX2_X1 port map( A => REGISTERS_12_41_port, B => n5833, S => n63, Z
                           => n3713);
   U4824 : MUX2_X1 port map( A => REGISTERS_12_40_port, B => n5834, S => n63, Z
                           => n3712);
   U4825 : MUX2_X1 port map( A => REGISTERS_12_39_port, B => n5835, S => n63, Z
                           => n3711);
   U4826 : MUX2_X1 port map( A => REGISTERS_12_38_port, B => n5836, S => n63, Z
                           => n3710);
   U4827 : MUX2_X1 port map( A => REGISTERS_12_37_port, B => n5837, S => n63, Z
                           => n3709);
   U4828 : MUX2_X1 port map( A => REGISTERS_12_36_port, B => n5838, S => n63, Z
                           => n3708);
   U4829 : MUX2_X1 port map( A => REGISTERS_12_35_port, B => n5839, S => n63, Z
                           => n3707);
   U4830 : MUX2_X1 port map( A => REGISTERS_12_34_port, B => n5840, S => n63, Z
                           => n3706);
   U4831 : MUX2_X1 port map( A => REGISTERS_12_33_port, B => n5841, S => n63, Z
                           => n3705);
   U4832 : MUX2_X1 port map( A => REGISTERS_12_32_port, B => n5842, S => n63, Z
                           => n3704);
   U4833 : MUX2_X1 port map( A => REGISTERS_12_31_port, B => n5843, S => n63, Z
                           => n3703);
   U4834 : MUX2_X1 port map( A => REGISTERS_12_30_port, B => n5844, S => n63, Z
                           => n3702);
   U4835 : MUX2_X1 port map( A => REGISTERS_12_29_port, B => n5845, S => n63, Z
                           => n3701);
   U4836 : MUX2_X1 port map( A => REGISTERS_12_28_port, B => n5846, S => n63, Z
                           => n3700);
   U4837 : MUX2_X1 port map( A => REGISTERS_12_27_port, B => n5847, S => n63, Z
                           => n3699);
   U4838 : MUX2_X1 port map( A => REGISTERS_12_26_port, B => n5848, S => n63, Z
                           => n3698);
   U4839 : MUX2_X1 port map( A => REGISTERS_12_25_port, B => n5849, S => n63, Z
                           => n3697);
   U4840 : MUX2_X1 port map( A => REGISTERS_12_24_port, B => n5850, S => n63, Z
                           => n3696);
   U4841 : MUX2_X1 port map( A => REGISTERS_12_23_port, B => n5851, S => n63, Z
                           => n3695);
   U4842 : MUX2_X1 port map( A => REGISTERS_12_22_port, B => n5852, S => n63, Z
                           => n3694);
   U4843 : MUX2_X1 port map( A => REGISTERS_12_21_port, B => n5853, S => n63, Z
                           => n3693);
   U4844 : MUX2_X1 port map( A => REGISTERS_12_20_port, B => n5854, S => n63, Z
                           => n3692);
   U4845 : MUX2_X1 port map( A => REGISTERS_12_19_port, B => n5855, S => n63, Z
                           => n3691);
   U4846 : MUX2_X1 port map( A => REGISTERS_12_18_port, B => n5856, S => n63, Z
                           => n3690);
   U4847 : MUX2_X1 port map( A => REGISTERS_12_17_port, B => n5857, S => n63, Z
                           => n3689);
   U4848 : MUX2_X1 port map( A => REGISTERS_12_16_port, B => n5858, S => n63, Z
                           => n3688);
   U4849 : MUX2_X1 port map( A => REGISTERS_12_15_port, B => n5859, S => n63, Z
                           => n3687);
   U4850 : MUX2_X1 port map( A => REGISTERS_12_14_port, B => n5860, S => n63, Z
                           => n3686);
   U4851 : MUX2_X1 port map( A => REGISTERS_12_13_port, B => n5861, S => n63, Z
                           => n3685);
   U4852 : MUX2_X1 port map( A => REGISTERS_12_12_port, B => n5862, S => n63, Z
                           => n3684);
   U4853 : MUX2_X1 port map( A => REGISTERS_12_11_port, B => n5863, S => n63, Z
                           => n3683);
   U4854 : MUX2_X1 port map( A => REGISTERS_12_10_port, B => n5864, S => n63, Z
                           => n3682);
   U4855 : MUX2_X1 port map( A => REGISTERS_12_9_port, B => n5865, S => n63, Z 
                           => n3681);
   U4856 : MUX2_X1 port map( A => REGISTERS_12_8_port, B => n5866, S => n63, Z 
                           => n3680);
   U4857 : MUX2_X1 port map( A => REGISTERS_12_7_port, B => n5867, S => n63, Z 
                           => n3679);
   U4858 : MUX2_X1 port map( A => REGISTERS_12_6_port, B => n5868, S => n63, Z 
                           => n3678);
   U4859 : MUX2_X1 port map( A => REGISTERS_12_5_port, B => n5869, S => n63, Z 
                           => n3677);
   U4860 : MUX2_X1 port map( A => REGISTERS_12_4_port, B => n5870, S => n63, Z 
                           => n3676);
   U4861 : MUX2_X1 port map( A => REGISTERS_12_3_port, B => n5871, S => n63, Z 
                           => n3675);
   U4862 : MUX2_X1 port map( A => REGISTERS_12_2_port, B => n5872, S => n63, Z 
                           => n3674);
   U4863 : MUX2_X1 port map( A => REGISTERS_12_1_port, B => n5873, S => n63, Z 
                           => n3673);
   U4864 : MUX2_X1 port map( A => REGISTERS_12_0_port, B => n5874, S => n63, Z 
                           => n3672);
   U4865 : OAI21_X1 port map( B1 => n5884, B2 => n5895, A => n5744, ZN => n5899
                           );
   U4866 : MUX2_X1 port map( A => REGISTERS_13_63_port, B => n5810, S => n65, Z
                           => n3671);
   U4867 : MUX2_X1 port map( A => REGISTERS_13_62_port, B => n5812, S => n65, Z
                           => n3670);
   U4868 : MUX2_X1 port map( A => REGISTERS_13_61_port, B => n5813, S => n65, Z
                           => n3669);
   U4869 : MUX2_X1 port map( A => REGISTERS_13_60_port, B => n5814, S => n65, Z
                           => n3668);
   U4870 : MUX2_X1 port map( A => REGISTERS_13_59_port, B => n5815, S => n65, Z
                           => n3667);
   U4871 : MUX2_X1 port map( A => REGISTERS_13_58_port, B => n5816, S => n65, Z
                           => n3666);
   U4872 : MUX2_X1 port map( A => REGISTERS_13_57_port, B => n5817, S => n65, Z
                           => n3665);
   U4873 : MUX2_X1 port map( A => REGISTERS_13_56_port, B => n5818, S => n65, Z
                           => n3664);
   U4874 : MUX2_X1 port map( A => REGISTERS_13_55_port, B => n5819, S => n65, Z
                           => n3663);
   U4875 : MUX2_X1 port map( A => REGISTERS_13_54_port, B => n5820, S => n65, Z
                           => n3662);
   U4876 : MUX2_X1 port map( A => REGISTERS_13_53_port, B => n5821, S => n65, Z
                           => n3661);
   U4877 : MUX2_X1 port map( A => REGISTERS_13_52_port, B => n5822, S => n65, Z
                           => n3660);
   U4878 : MUX2_X1 port map( A => REGISTERS_13_51_port, B => n5823, S => n65, Z
                           => n3659);
   U4879 : MUX2_X1 port map( A => REGISTERS_13_50_port, B => n5824, S => n65, Z
                           => n3658);
   U4880 : MUX2_X1 port map( A => REGISTERS_13_49_port, B => n5825, S => n65, Z
                           => n3657);
   U4881 : MUX2_X1 port map( A => REGISTERS_13_48_port, B => n5826, S => n65, Z
                           => n3656);
   U4882 : MUX2_X1 port map( A => REGISTERS_13_47_port, B => n5827, S => n65, Z
                           => n3655);
   U4883 : MUX2_X1 port map( A => REGISTERS_13_46_port, B => n5828, S => n65, Z
                           => n3654);
   U4884 : MUX2_X1 port map( A => REGISTERS_13_45_port, B => n5829, S => n65, Z
                           => n3653);
   U4885 : MUX2_X1 port map( A => REGISTERS_13_44_port, B => n5830, S => n65, Z
                           => n3652);
   U4886 : MUX2_X1 port map( A => REGISTERS_13_43_port, B => n5831, S => n65, Z
                           => n3651);
   U4887 : MUX2_X1 port map( A => REGISTERS_13_42_port, B => n5832, S => n65, Z
                           => n3650);
   U4888 : MUX2_X1 port map( A => REGISTERS_13_41_port, B => n5833, S => n65, Z
                           => n3649);
   U4889 : MUX2_X1 port map( A => REGISTERS_13_40_port, B => n5834, S => n65, Z
                           => n3648);
   U4890 : MUX2_X1 port map( A => REGISTERS_13_39_port, B => n5835, S => n65, Z
                           => n3647);
   U4891 : MUX2_X1 port map( A => REGISTERS_13_38_port, B => n5836, S => n65, Z
                           => n3646);
   U4892 : MUX2_X1 port map( A => REGISTERS_13_37_port, B => n5837, S => n65, Z
                           => n3645);
   U4893 : MUX2_X1 port map( A => REGISTERS_13_36_port, B => n5838, S => n65, Z
                           => n3644);
   U4894 : MUX2_X1 port map( A => REGISTERS_13_35_port, B => n5839, S => n65, Z
                           => n3643);
   U4895 : MUX2_X1 port map( A => REGISTERS_13_34_port, B => n5840, S => n65, Z
                           => n3642);
   U4896 : MUX2_X1 port map( A => REGISTERS_13_33_port, B => n5841, S => n65, Z
                           => n3641);
   U4897 : MUX2_X1 port map( A => REGISTERS_13_32_port, B => n5842, S => n65, Z
                           => n3640);
   U4898 : MUX2_X1 port map( A => REGISTERS_13_31_port, B => n5843, S => n65, Z
                           => n3639);
   U4899 : MUX2_X1 port map( A => REGISTERS_13_30_port, B => n5844, S => n65, Z
                           => n3638);
   U4900 : MUX2_X1 port map( A => REGISTERS_13_29_port, B => n5845, S => n65, Z
                           => n3637);
   U4901 : MUX2_X1 port map( A => REGISTERS_13_28_port, B => n5846, S => n65, Z
                           => n3636);
   U4902 : MUX2_X1 port map( A => REGISTERS_13_27_port, B => n5847, S => n65, Z
                           => n3635);
   U4903 : MUX2_X1 port map( A => REGISTERS_13_26_port, B => n5848, S => n65, Z
                           => n3634);
   U4904 : MUX2_X1 port map( A => REGISTERS_13_25_port, B => n5849, S => n65, Z
                           => n3633);
   U4905 : MUX2_X1 port map( A => REGISTERS_13_24_port, B => n5850, S => n65, Z
                           => n3632);
   U4906 : MUX2_X1 port map( A => REGISTERS_13_23_port, B => n5851, S => n65, Z
                           => n3631);
   U4907 : MUX2_X1 port map( A => REGISTERS_13_22_port, B => n5852, S => n65, Z
                           => n3630);
   U4908 : MUX2_X1 port map( A => REGISTERS_13_21_port, B => n5853, S => n65, Z
                           => n3629);
   U4909 : MUX2_X1 port map( A => REGISTERS_13_20_port, B => n5854, S => n65, Z
                           => n3628);
   U4910 : MUX2_X1 port map( A => REGISTERS_13_19_port, B => n5855, S => n65, Z
                           => n3627);
   U4911 : MUX2_X1 port map( A => REGISTERS_13_18_port, B => n5856, S => n65, Z
                           => n3626);
   U4912 : MUX2_X1 port map( A => REGISTERS_13_17_port, B => n5857, S => n65, Z
                           => n3625);
   U4913 : MUX2_X1 port map( A => REGISTERS_13_16_port, B => n5858, S => n65, Z
                           => n3624);
   U4914 : MUX2_X1 port map( A => REGISTERS_13_15_port, B => n5859, S => n65, Z
                           => n3623);
   U4915 : MUX2_X1 port map( A => REGISTERS_13_14_port, B => n5860, S => n65, Z
                           => n3622);
   U4916 : MUX2_X1 port map( A => REGISTERS_13_13_port, B => n5861, S => n65, Z
                           => n3621);
   U4917 : MUX2_X1 port map( A => REGISTERS_13_12_port, B => n5862, S => n65, Z
                           => n3620);
   U4918 : MUX2_X1 port map( A => REGISTERS_13_11_port, B => n5863, S => n65, Z
                           => n3619);
   U4919 : MUX2_X1 port map( A => REGISTERS_13_10_port, B => n5864, S => n65, Z
                           => n3618);
   U4920 : MUX2_X1 port map( A => REGISTERS_13_9_port, B => n5865, S => n65, Z 
                           => n3617);
   U4921 : MUX2_X1 port map( A => REGISTERS_13_8_port, B => n5866, S => n65, Z 
                           => n3616);
   U4922 : MUX2_X1 port map( A => REGISTERS_13_7_port, B => n5867, S => n65, Z 
                           => n3615);
   U4923 : MUX2_X1 port map( A => REGISTERS_13_6_port, B => n5868, S => n65, Z 
                           => n3614);
   U4924 : MUX2_X1 port map( A => REGISTERS_13_5_port, B => n5869, S => n65, Z 
                           => n3613);
   U4925 : MUX2_X1 port map( A => REGISTERS_13_4_port, B => n5870, S => n65, Z 
                           => n3612);
   U4926 : MUX2_X1 port map( A => REGISTERS_13_3_port, B => n5871, S => n65, Z 
                           => n3611);
   U4927 : MUX2_X1 port map( A => REGISTERS_13_2_port, B => n5872, S => n65, Z 
                           => n3610);
   U4928 : MUX2_X1 port map( A => REGISTERS_13_1_port, B => n5873, S => n65, Z 
                           => n3609);
   U4929 : MUX2_X1 port map( A => REGISTERS_13_0_port, B => n5874, S => n65, Z 
                           => n3608);
   U4930 : OAI21_X1 port map( B1 => n5886, B2 => n5895, A => n5744, ZN => n5900
                           );
   U4931 : MUX2_X1 port map( A => REGISTERS_14_63_port, B => n5810, S => n67, Z
                           => n3607);
   U4932 : MUX2_X1 port map( A => REGISTERS_14_62_port, B => n5812, S => n67, Z
                           => n3606);
   U4933 : MUX2_X1 port map( A => REGISTERS_14_61_port, B => n5813, S => n67, Z
                           => n3605);
   U4934 : MUX2_X1 port map( A => REGISTERS_14_60_port, B => n5814, S => n67, Z
                           => n3604);
   U4935 : MUX2_X1 port map( A => REGISTERS_14_59_port, B => n5815, S => n67, Z
                           => n3603);
   U4936 : MUX2_X1 port map( A => REGISTERS_14_58_port, B => n5816, S => n67, Z
                           => n3602);
   U4937 : MUX2_X1 port map( A => REGISTERS_14_57_port, B => n5817, S => n67, Z
                           => n3601);
   U4938 : MUX2_X1 port map( A => REGISTERS_14_56_port, B => n5818, S => n67, Z
                           => n3600);
   U4939 : MUX2_X1 port map( A => REGISTERS_14_55_port, B => n5819, S => n67, Z
                           => n3599);
   U4940 : MUX2_X1 port map( A => REGISTERS_14_54_port, B => n5820, S => n67, Z
                           => n3598);
   U4941 : MUX2_X1 port map( A => REGISTERS_14_53_port, B => n5821, S => n67, Z
                           => n3597);
   U4942 : MUX2_X1 port map( A => REGISTERS_14_52_port, B => n5822, S => n67, Z
                           => n3596);
   U4943 : MUX2_X1 port map( A => REGISTERS_14_51_port, B => n5823, S => n67, Z
                           => n3595);
   U4944 : MUX2_X1 port map( A => REGISTERS_14_50_port, B => n5824, S => n67, Z
                           => n3594);
   U4945 : MUX2_X1 port map( A => REGISTERS_14_49_port, B => n5825, S => n67, Z
                           => n3593);
   U4946 : MUX2_X1 port map( A => REGISTERS_14_48_port, B => n5826, S => n67, Z
                           => n3592);
   U4947 : MUX2_X1 port map( A => REGISTERS_14_47_port, B => n5827, S => n67, Z
                           => n3591);
   U4948 : MUX2_X1 port map( A => REGISTERS_14_46_port, B => n5828, S => n67, Z
                           => n3590);
   U4949 : MUX2_X1 port map( A => REGISTERS_14_45_port, B => n5829, S => n67, Z
                           => n3589);
   U4950 : MUX2_X1 port map( A => REGISTERS_14_44_port, B => n5830, S => n67, Z
                           => n3588);
   U4951 : MUX2_X1 port map( A => REGISTERS_14_43_port, B => n5831, S => n67, Z
                           => n3587);
   U4952 : MUX2_X1 port map( A => REGISTERS_14_42_port, B => n5832, S => n67, Z
                           => n3586);
   U4953 : MUX2_X1 port map( A => REGISTERS_14_41_port, B => n5833, S => n67, Z
                           => n3585);
   U4954 : MUX2_X1 port map( A => REGISTERS_14_40_port, B => n5834, S => n67, Z
                           => n3584);
   U4955 : MUX2_X1 port map( A => REGISTERS_14_39_port, B => n5835, S => n67, Z
                           => n3583);
   U4956 : MUX2_X1 port map( A => REGISTERS_14_38_port, B => n5836, S => n67, Z
                           => n3582);
   U4957 : MUX2_X1 port map( A => REGISTERS_14_37_port, B => n5837, S => n67, Z
                           => n3581);
   U4958 : MUX2_X1 port map( A => REGISTERS_14_36_port, B => n5838, S => n67, Z
                           => n3580);
   U4959 : MUX2_X1 port map( A => REGISTERS_14_35_port, B => n5839, S => n67, Z
                           => n3579);
   U4960 : MUX2_X1 port map( A => REGISTERS_14_34_port, B => n5840, S => n67, Z
                           => n3578);
   U4961 : MUX2_X1 port map( A => REGISTERS_14_33_port, B => n5841, S => n67, Z
                           => n3577);
   U4962 : MUX2_X1 port map( A => REGISTERS_14_32_port, B => n5842, S => n67, Z
                           => n3576);
   U4963 : MUX2_X1 port map( A => REGISTERS_14_31_port, B => n5843, S => n67, Z
                           => n3575);
   U4964 : MUX2_X1 port map( A => REGISTERS_14_30_port, B => n5844, S => n67, Z
                           => n3574);
   U4965 : MUX2_X1 port map( A => REGISTERS_14_29_port, B => n5845, S => n67, Z
                           => n3573);
   U4966 : MUX2_X1 port map( A => REGISTERS_14_28_port, B => n5846, S => n67, Z
                           => n3572);
   U4967 : MUX2_X1 port map( A => REGISTERS_14_27_port, B => n5847, S => n67, Z
                           => n3571);
   U4968 : MUX2_X1 port map( A => REGISTERS_14_26_port, B => n5848, S => n67, Z
                           => n3570);
   U4969 : MUX2_X1 port map( A => REGISTERS_14_25_port, B => n5849, S => n67, Z
                           => n3569);
   U4970 : MUX2_X1 port map( A => REGISTERS_14_24_port, B => n5850, S => n67, Z
                           => n3568);
   U4971 : MUX2_X1 port map( A => REGISTERS_14_23_port, B => n5851, S => n67, Z
                           => n3567);
   U4972 : MUX2_X1 port map( A => REGISTERS_14_22_port, B => n5852, S => n67, Z
                           => n3566);
   U4973 : MUX2_X1 port map( A => REGISTERS_14_21_port, B => n5853, S => n67, Z
                           => n3565);
   U4974 : MUX2_X1 port map( A => REGISTERS_14_20_port, B => n5854, S => n67, Z
                           => n3564);
   U4975 : MUX2_X1 port map( A => REGISTERS_14_19_port, B => n5855, S => n67, Z
                           => n3563);
   U4976 : MUX2_X1 port map( A => REGISTERS_14_18_port, B => n5856, S => n67, Z
                           => n3562);
   U4977 : MUX2_X1 port map( A => REGISTERS_14_17_port, B => n5857, S => n67, Z
                           => n3561);
   U4978 : MUX2_X1 port map( A => REGISTERS_14_16_port, B => n5858, S => n67, Z
                           => n3560);
   U4979 : MUX2_X1 port map( A => REGISTERS_14_15_port, B => n5859, S => n67, Z
                           => n3559);
   U4980 : MUX2_X1 port map( A => REGISTERS_14_14_port, B => n5860, S => n67, Z
                           => n3558);
   U4981 : MUX2_X1 port map( A => REGISTERS_14_13_port, B => n5861, S => n67, Z
                           => n3557);
   U4982 : MUX2_X1 port map( A => REGISTERS_14_12_port, B => n5862, S => n67, Z
                           => n3556);
   U4983 : MUX2_X1 port map( A => REGISTERS_14_11_port, B => n5863, S => n67, Z
                           => n3555);
   U4984 : MUX2_X1 port map( A => REGISTERS_14_10_port, B => n5864, S => n67, Z
                           => n3554);
   U4985 : MUX2_X1 port map( A => REGISTERS_14_9_port, B => n5865, S => n67, Z 
                           => n3553);
   U4986 : MUX2_X1 port map( A => REGISTERS_14_8_port, B => n5866, S => n67, Z 
                           => n3552);
   U4987 : MUX2_X1 port map( A => REGISTERS_14_7_port, B => n5867, S => n67, Z 
                           => n3551);
   U4988 : MUX2_X1 port map( A => REGISTERS_14_6_port, B => n5868, S => n67, Z 
                           => n3550);
   U4989 : MUX2_X1 port map( A => REGISTERS_14_5_port, B => n5869, S => n67, Z 
                           => n3549);
   U4990 : MUX2_X1 port map( A => REGISTERS_14_4_port, B => n5870, S => n67, Z 
                           => n3548);
   U4991 : MUX2_X1 port map( A => REGISTERS_14_3_port, B => n5871, S => n67, Z 
                           => n3547);
   U4992 : MUX2_X1 port map( A => REGISTERS_14_2_port, B => n5872, S => n67, Z 
                           => n3546);
   U4993 : MUX2_X1 port map( A => REGISTERS_14_1_port, B => n5873, S => n67, Z 
                           => n3545);
   U4994 : MUX2_X1 port map( A => REGISTERS_14_0_port, B => n5874, S => n67, Z 
                           => n3544);
   U4995 : OAI21_X1 port map( B1 => n5888, B2 => n5895, A => n5744, ZN => n5901
                           );
   U4996 : MUX2_X1 port map( A => REGISTERS_15_63_port, B => n5810, S => n53, Z
                           => n3543);
   U4997 : MUX2_X1 port map( A => REGISTERS_15_62_port, B => n5812, S => n53, Z
                           => n3542);
   U4998 : MUX2_X1 port map( A => REGISTERS_15_61_port, B => n5813, S => n53, Z
                           => n3541);
   U4999 : MUX2_X1 port map( A => REGISTERS_15_60_port, B => n5814, S => n53, Z
                           => n3540);
   U5000 : MUX2_X1 port map( A => REGISTERS_15_59_port, B => n5815, S => n53, Z
                           => n3539);
   U5001 : MUX2_X1 port map( A => REGISTERS_15_58_port, B => n5816, S => n53, Z
                           => n3538);
   U5002 : MUX2_X1 port map( A => REGISTERS_15_57_port, B => n5817, S => n53, Z
                           => n3537);
   U5003 : MUX2_X1 port map( A => REGISTERS_15_56_port, B => n5818, S => n53, Z
                           => n3536);
   U5004 : MUX2_X1 port map( A => REGISTERS_15_55_port, B => n5819, S => n53, Z
                           => n3535);
   U5005 : MUX2_X1 port map( A => REGISTERS_15_54_port, B => n5820, S => n53, Z
                           => n3534);
   U5006 : MUX2_X1 port map( A => REGISTERS_15_53_port, B => n5821, S => n53, Z
                           => n3533);
   U5007 : MUX2_X1 port map( A => REGISTERS_15_52_port, B => n5822, S => n53, Z
                           => n3532);
   U5008 : MUX2_X1 port map( A => REGISTERS_15_51_port, B => n5823, S => n53, Z
                           => n3531);
   U5009 : MUX2_X1 port map( A => REGISTERS_15_50_port, B => n5824, S => n53, Z
                           => n3530);
   U5010 : MUX2_X1 port map( A => REGISTERS_15_49_port, B => n5825, S => n53, Z
                           => n3529);
   U5011 : MUX2_X1 port map( A => REGISTERS_15_48_port, B => n5826, S => n53, Z
                           => n3528);
   U5012 : MUX2_X1 port map( A => REGISTERS_15_47_port, B => n5827, S => n53, Z
                           => n3527);
   U5013 : MUX2_X1 port map( A => REGISTERS_15_46_port, B => n5828, S => n53, Z
                           => n3526);
   U5014 : MUX2_X1 port map( A => REGISTERS_15_45_port, B => n5829, S => n53, Z
                           => n3525);
   U5015 : MUX2_X1 port map( A => REGISTERS_15_44_port, B => n5830, S => n53, Z
                           => n3524);
   U5016 : MUX2_X1 port map( A => REGISTERS_15_43_port, B => n5831, S => n53, Z
                           => n3523);
   U5017 : MUX2_X1 port map( A => REGISTERS_15_42_port, B => n5832, S => n53, Z
                           => n3522);
   U5018 : MUX2_X1 port map( A => REGISTERS_15_41_port, B => n5833, S => n53, Z
                           => n3521);
   U5019 : MUX2_X1 port map( A => REGISTERS_15_40_port, B => n5834, S => n53, Z
                           => n3520);
   U5020 : MUX2_X1 port map( A => REGISTERS_15_39_port, B => n5835, S => n53, Z
                           => n3519);
   U5021 : MUX2_X1 port map( A => REGISTERS_15_38_port, B => n5836, S => n53, Z
                           => n3518);
   U5022 : MUX2_X1 port map( A => REGISTERS_15_37_port, B => n5837, S => n53, Z
                           => n3517);
   U5023 : MUX2_X1 port map( A => REGISTERS_15_36_port, B => n5838, S => n53, Z
                           => n3516);
   U5024 : MUX2_X1 port map( A => REGISTERS_15_35_port, B => n5839, S => n53, Z
                           => n3515);
   U5025 : MUX2_X1 port map( A => REGISTERS_15_34_port, B => n5840, S => n53, Z
                           => n3514);
   U5026 : MUX2_X1 port map( A => REGISTERS_15_33_port, B => n5841, S => n53, Z
                           => n3513);
   U5027 : MUX2_X1 port map( A => REGISTERS_15_32_port, B => n5842, S => n53, Z
                           => n3512);
   U5028 : MUX2_X1 port map( A => REGISTERS_15_31_port, B => n5843, S => n53, Z
                           => n3511);
   U5029 : MUX2_X1 port map( A => REGISTERS_15_30_port, B => n5844, S => n53, Z
                           => n3510);
   U5030 : MUX2_X1 port map( A => REGISTERS_15_29_port, B => n5845, S => n53, Z
                           => n3509);
   U5031 : MUX2_X1 port map( A => REGISTERS_15_28_port, B => n5846, S => n53, Z
                           => n3508);
   U5032 : MUX2_X1 port map( A => REGISTERS_15_27_port, B => n5847, S => n53, Z
                           => n3507);
   U5033 : MUX2_X1 port map( A => REGISTERS_15_26_port, B => n5848, S => n53, Z
                           => n3506);
   U5034 : MUX2_X1 port map( A => REGISTERS_15_25_port, B => n5849, S => n53, Z
                           => n3505);
   U5035 : MUX2_X1 port map( A => REGISTERS_15_24_port, B => n5850, S => n53, Z
                           => n3504);
   U5036 : MUX2_X1 port map( A => REGISTERS_15_23_port, B => n5851, S => n53, Z
                           => n3503);
   U5037 : MUX2_X1 port map( A => REGISTERS_15_22_port, B => n5852, S => n53, Z
                           => n3502);
   U5038 : MUX2_X1 port map( A => REGISTERS_15_21_port, B => n5853, S => n53, Z
                           => n3501);
   U5039 : MUX2_X1 port map( A => REGISTERS_15_20_port, B => n5854, S => n53, Z
                           => n3500);
   U5040 : MUX2_X1 port map( A => REGISTERS_15_19_port, B => n5855, S => n53, Z
                           => n3499);
   U5041 : MUX2_X1 port map( A => REGISTERS_15_18_port, B => n5856, S => n53, Z
                           => n3498);
   U5042 : MUX2_X1 port map( A => REGISTERS_15_17_port, B => n5857, S => n53, Z
                           => n3497);
   U5043 : MUX2_X1 port map( A => REGISTERS_15_16_port, B => n5858, S => n53, Z
                           => n3496);
   U5044 : MUX2_X1 port map( A => REGISTERS_15_15_port, B => n5859, S => n53, Z
                           => n3495);
   U5045 : MUX2_X1 port map( A => REGISTERS_15_14_port, B => n5860, S => n53, Z
                           => n3494);
   U5046 : MUX2_X1 port map( A => REGISTERS_15_13_port, B => n5861, S => n53, Z
                           => n3493);
   U5047 : MUX2_X1 port map( A => REGISTERS_15_12_port, B => n5862, S => n53, Z
                           => n3492);
   U5048 : MUX2_X1 port map( A => REGISTERS_15_11_port, B => n5863, S => n53, Z
                           => n3491);
   U5049 : MUX2_X1 port map( A => REGISTERS_15_10_port, B => n5864, S => n53, Z
                           => n3490);
   U5050 : MUX2_X1 port map( A => REGISTERS_15_9_port, B => n5865, S => n53, Z 
                           => n3489);
   U5051 : MUX2_X1 port map( A => REGISTERS_15_8_port, B => n5866, S => n53, Z 
                           => n3488);
   U5052 : MUX2_X1 port map( A => REGISTERS_15_7_port, B => n5867, S => n53, Z 
                           => n3487);
   U5053 : MUX2_X1 port map( A => REGISTERS_15_6_port, B => n5868, S => n53, Z 
                           => n3486);
   U5054 : MUX2_X1 port map( A => REGISTERS_15_5_port, B => n5869, S => n53, Z 
                           => n3485);
   U5055 : MUX2_X1 port map( A => REGISTERS_15_4_port, B => n5870, S => n53, Z 
                           => n3484);
   U5056 : MUX2_X1 port map( A => REGISTERS_15_3_port, B => n5871, S => n53, Z 
                           => n3483);
   U5057 : MUX2_X1 port map( A => REGISTERS_15_2_port, B => n5872, S => n53, Z 
                           => n3482);
   U5058 : MUX2_X1 port map( A => REGISTERS_15_1_port, B => n5873, S => n53, Z 
                           => n3481);
   U5059 : MUX2_X1 port map( A => REGISTERS_15_0_port, B => n5874, S => n53, Z 
                           => n3480);
   U5060 : OAI21_X1 port map( B1 => n5890, B2 => n5895, A => n5744, ZN => n5902
                           );
   U5061 : NAND3_X1 port map( A1 => n5893, A2 => n5892, A3 => ADD_WR(3), ZN => 
                           n5895);
   U5062 : INV_X1 port map( A => ADD_WR(4), ZN => n5892);
   U5063 : MUX2_X1 port map( A => REGISTERS_16_63_port, B => n5810, S => n55, Z
                           => n3479);
   U5064 : MUX2_X1 port map( A => REGISTERS_16_62_port, B => n5812, S => n55, Z
                           => n3478);
   U5065 : MUX2_X1 port map( A => REGISTERS_16_61_port, B => n5813, S => n55, Z
                           => n3477);
   U5066 : MUX2_X1 port map( A => REGISTERS_16_60_port, B => n5814, S => n55, Z
                           => n3476);
   U5067 : MUX2_X1 port map( A => REGISTERS_16_59_port, B => n5815, S => n55, Z
                           => n3475);
   U5068 : MUX2_X1 port map( A => REGISTERS_16_58_port, B => n5816, S => n55, Z
                           => n3474);
   U5069 : MUX2_X1 port map( A => REGISTERS_16_57_port, B => n5817, S => n55, Z
                           => n3473);
   U5070 : MUX2_X1 port map( A => REGISTERS_16_56_port, B => n5818, S => n55, Z
                           => n3472);
   U5071 : MUX2_X1 port map( A => REGISTERS_16_55_port, B => n5819, S => n55, Z
                           => n3471);
   U5072 : MUX2_X1 port map( A => REGISTERS_16_54_port, B => n5820, S => n55, Z
                           => n3470);
   U5073 : MUX2_X1 port map( A => REGISTERS_16_53_port, B => n5821, S => n55, Z
                           => n3469);
   U5074 : MUX2_X1 port map( A => REGISTERS_16_52_port, B => n5822, S => n55, Z
                           => n3468);
   U5075 : MUX2_X1 port map( A => REGISTERS_16_51_port, B => n5823, S => n55, Z
                           => n3467);
   U5076 : MUX2_X1 port map( A => REGISTERS_16_50_port, B => n5824, S => n55, Z
                           => n3466);
   U5077 : MUX2_X1 port map( A => REGISTERS_16_49_port, B => n5825, S => n55, Z
                           => n3465);
   U5078 : MUX2_X1 port map( A => REGISTERS_16_48_port, B => n5826, S => n55, Z
                           => n3464);
   U5079 : MUX2_X1 port map( A => REGISTERS_16_47_port, B => n5827, S => n55, Z
                           => n3463);
   U5080 : MUX2_X1 port map( A => REGISTERS_16_46_port, B => n5828, S => n55, Z
                           => n3462);
   U5081 : MUX2_X1 port map( A => REGISTERS_16_45_port, B => n5829, S => n55, Z
                           => n3461);
   U5082 : MUX2_X1 port map( A => REGISTERS_16_44_port, B => n5830, S => n55, Z
                           => n3460);
   U5083 : MUX2_X1 port map( A => REGISTERS_16_43_port, B => n5831, S => n55, Z
                           => n3459);
   U5084 : MUX2_X1 port map( A => REGISTERS_16_42_port, B => n5832, S => n55, Z
                           => n3458);
   U5085 : MUX2_X1 port map( A => REGISTERS_16_41_port, B => n5833, S => n55, Z
                           => n3457);
   U5086 : MUX2_X1 port map( A => REGISTERS_16_40_port, B => n5834, S => n55, Z
                           => n3456);
   U5087 : MUX2_X1 port map( A => REGISTERS_16_39_port, B => n5835, S => n55, Z
                           => n3455);
   U5088 : MUX2_X1 port map( A => REGISTERS_16_38_port, B => n5836, S => n55, Z
                           => n3454);
   U5089 : MUX2_X1 port map( A => REGISTERS_16_37_port, B => n5837, S => n55, Z
                           => n3453);
   U5090 : MUX2_X1 port map( A => REGISTERS_16_36_port, B => n5838, S => n55, Z
                           => n3452);
   U5091 : MUX2_X1 port map( A => REGISTERS_16_35_port, B => n5839, S => n55, Z
                           => n3451);
   U5092 : MUX2_X1 port map( A => REGISTERS_16_34_port, B => n5840, S => n55, Z
                           => n3450);
   U5093 : MUX2_X1 port map( A => REGISTERS_16_33_port, B => n5841, S => n55, Z
                           => n3449);
   U5094 : MUX2_X1 port map( A => REGISTERS_16_32_port, B => n5842, S => n55, Z
                           => n3448);
   U5095 : MUX2_X1 port map( A => REGISTERS_16_31_port, B => n5843, S => n55, Z
                           => n3447);
   U5096 : MUX2_X1 port map( A => REGISTERS_16_30_port, B => n5844, S => n55, Z
                           => n3446);
   U5097 : MUX2_X1 port map( A => REGISTERS_16_29_port, B => n5845, S => n55, Z
                           => n3445);
   U5098 : MUX2_X1 port map( A => REGISTERS_16_28_port, B => n5846, S => n55, Z
                           => n3444);
   U5099 : MUX2_X1 port map( A => REGISTERS_16_27_port, B => n5847, S => n55, Z
                           => n3443);
   U5100 : MUX2_X1 port map( A => REGISTERS_16_26_port, B => n5848, S => n55, Z
                           => n3442);
   U5101 : MUX2_X1 port map( A => REGISTERS_16_25_port, B => n5849, S => n55, Z
                           => n3441);
   U5102 : MUX2_X1 port map( A => REGISTERS_16_24_port, B => n5850, S => n55, Z
                           => n3440);
   U5103 : MUX2_X1 port map( A => REGISTERS_16_23_port, B => n5851, S => n55, Z
                           => n3439);
   U5104 : MUX2_X1 port map( A => REGISTERS_16_22_port, B => n5852, S => n55, Z
                           => n3438);
   U5105 : MUX2_X1 port map( A => REGISTERS_16_21_port, B => n5853, S => n55, Z
                           => n3437);
   U5106 : MUX2_X1 port map( A => REGISTERS_16_20_port, B => n5854, S => n55, Z
                           => n3436);
   U5107 : MUX2_X1 port map( A => REGISTERS_16_19_port, B => n5855, S => n55, Z
                           => n3435);
   U5108 : MUX2_X1 port map( A => REGISTERS_16_18_port, B => n5856, S => n55, Z
                           => n3434);
   U5109 : MUX2_X1 port map( A => REGISTERS_16_17_port, B => n5857, S => n55, Z
                           => n3433);
   U5110 : MUX2_X1 port map( A => REGISTERS_16_16_port, B => n5858, S => n55, Z
                           => n3432);
   U5111 : MUX2_X1 port map( A => REGISTERS_16_15_port, B => n5859, S => n55, Z
                           => n3431);
   U5112 : MUX2_X1 port map( A => REGISTERS_16_14_port, B => n5860, S => n55, Z
                           => n3430);
   U5113 : MUX2_X1 port map( A => REGISTERS_16_13_port, B => n5861, S => n55, Z
                           => n3429);
   U5114 : MUX2_X1 port map( A => REGISTERS_16_12_port, B => n5862, S => n55, Z
                           => n3428);
   U5115 : MUX2_X1 port map( A => REGISTERS_16_11_port, B => n5863, S => n55, Z
                           => n3427);
   U5116 : MUX2_X1 port map( A => REGISTERS_16_10_port, B => n5864, S => n55, Z
                           => n3426);
   U5117 : MUX2_X1 port map( A => REGISTERS_16_9_port, B => n5865, S => n55, Z 
                           => n3425);
   U5118 : MUX2_X1 port map( A => REGISTERS_16_8_port, B => n5866, S => n55, Z 
                           => n3424);
   U5119 : MUX2_X1 port map( A => REGISTERS_16_7_port, B => n5867, S => n55, Z 
                           => n3423);
   U5120 : MUX2_X1 port map( A => REGISTERS_16_6_port, B => n5868, S => n55, Z 
                           => n3422);
   U5121 : MUX2_X1 port map( A => REGISTERS_16_5_port, B => n5869, S => n55, Z 
                           => n3421);
   U5122 : MUX2_X1 port map( A => REGISTERS_16_4_port, B => n5870, S => n55, Z 
                           => n3420);
   U5123 : MUX2_X1 port map( A => REGISTERS_16_3_port, B => n5871, S => n55, Z 
                           => n3419);
   U5124 : MUX2_X1 port map( A => REGISTERS_16_2_port, B => n5872, S => n55, Z 
                           => n3418);
   U5125 : MUX2_X1 port map( A => REGISTERS_16_1_port, B => n5873, S => n55, Z 
                           => n3417);
   U5126 : MUX2_X1 port map( A => REGISTERS_16_0_port, B => n5874, S => n55, Z 
                           => n3416);
   U5127 : OAI21_X1 port map( B1 => n5876, B2 => n5904, A => n5744, ZN => n5903
                           );
   U5128 : MUX2_X1 port map( A => REGISTERS_17_63_port, B => n5810, S => n57, Z
                           => n3415);
   U5129 : MUX2_X1 port map( A => REGISTERS_17_62_port, B => n5812, S => n57, Z
                           => n3414);
   U5130 : MUX2_X1 port map( A => REGISTERS_17_61_port, B => n5813, S => n57, Z
                           => n3413);
   U5131 : MUX2_X1 port map( A => REGISTERS_17_60_port, B => n5814, S => n57, Z
                           => n3412);
   U5132 : MUX2_X1 port map( A => REGISTERS_17_59_port, B => n5815, S => n57, Z
                           => n3411);
   U5133 : MUX2_X1 port map( A => REGISTERS_17_58_port, B => n5816, S => n57, Z
                           => n3410);
   U5134 : MUX2_X1 port map( A => REGISTERS_17_57_port, B => n5817, S => n57, Z
                           => n3409);
   U5135 : MUX2_X1 port map( A => REGISTERS_17_56_port, B => n5818, S => n57, Z
                           => n3408);
   U5136 : MUX2_X1 port map( A => REGISTERS_17_55_port, B => n5819, S => n57, Z
                           => n3407);
   U5137 : MUX2_X1 port map( A => REGISTERS_17_54_port, B => n5820, S => n57, Z
                           => n3406);
   U5138 : MUX2_X1 port map( A => REGISTERS_17_53_port, B => n5821, S => n57, Z
                           => n3405);
   U5139 : MUX2_X1 port map( A => REGISTERS_17_52_port, B => n5822, S => n57, Z
                           => n3404);
   U5140 : MUX2_X1 port map( A => REGISTERS_17_51_port, B => n5823, S => n57, Z
                           => n3403);
   U5141 : MUX2_X1 port map( A => REGISTERS_17_50_port, B => n5824, S => n57, Z
                           => n3402);
   U5142 : MUX2_X1 port map( A => REGISTERS_17_49_port, B => n5825, S => n57, Z
                           => n3401);
   U5143 : MUX2_X1 port map( A => REGISTERS_17_48_port, B => n5826, S => n57, Z
                           => n3400);
   U5144 : MUX2_X1 port map( A => REGISTERS_17_47_port, B => n5827, S => n57, Z
                           => n3399);
   U5145 : MUX2_X1 port map( A => REGISTERS_17_46_port, B => n5828, S => n57, Z
                           => n3398);
   U5146 : MUX2_X1 port map( A => REGISTERS_17_45_port, B => n5829, S => n57, Z
                           => n3397);
   U5147 : MUX2_X1 port map( A => REGISTERS_17_44_port, B => n5830, S => n57, Z
                           => n3396);
   U5148 : MUX2_X1 port map( A => REGISTERS_17_43_port, B => n5831, S => n57, Z
                           => n3395);
   U5149 : MUX2_X1 port map( A => REGISTERS_17_42_port, B => n5832, S => n57, Z
                           => n3394);
   U5150 : MUX2_X1 port map( A => REGISTERS_17_41_port, B => n5833, S => n57, Z
                           => n3393);
   U5151 : MUX2_X1 port map( A => REGISTERS_17_40_port, B => n5834, S => n57, Z
                           => n3392);
   U5152 : MUX2_X1 port map( A => REGISTERS_17_39_port, B => n5835, S => n57, Z
                           => n3391);
   U5153 : MUX2_X1 port map( A => REGISTERS_17_38_port, B => n5836, S => n57, Z
                           => n3390);
   U5154 : MUX2_X1 port map( A => REGISTERS_17_37_port, B => n5837, S => n57, Z
                           => n3389);
   U5155 : MUX2_X1 port map( A => REGISTERS_17_36_port, B => n5838, S => n57, Z
                           => n3388);
   U5156 : MUX2_X1 port map( A => REGISTERS_17_35_port, B => n5839, S => n57, Z
                           => n3387);
   U5157 : MUX2_X1 port map( A => REGISTERS_17_34_port, B => n5840, S => n57, Z
                           => n3386);
   U5158 : MUX2_X1 port map( A => REGISTERS_17_33_port, B => n5841, S => n57, Z
                           => n3385);
   U5159 : MUX2_X1 port map( A => REGISTERS_17_32_port, B => n5842, S => n57, Z
                           => n3384);
   U5160 : MUX2_X1 port map( A => REGISTERS_17_31_port, B => n5843, S => n57, Z
                           => n3383);
   U5161 : MUX2_X1 port map( A => REGISTERS_17_30_port, B => n5844, S => n57, Z
                           => n3382);
   U5162 : MUX2_X1 port map( A => REGISTERS_17_29_port, B => n5845, S => n57, Z
                           => n3381);
   U5163 : MUX2_X1 port map( A => REGISTERS_17_28_port, B => n5846, S => n57, Z
                           => n3380);
   U5164 : MUX2_X1 port map( A => REGISTERS_17_27_port, B => n5847, S => n57, Z
                           => n3379);
   U5165 : MUX2_X1 port map( A => REGISTERS_17_26_port, B => n5848, S => n57, Z
                           => n3378);
   U5166 : MUX2_X1 port map( A => REGISTERS_17_25_port, B => n5849, S => n57, Z
                           => n3377);
   U5167 : MUX2_X1 port map( A => REGISTERS_17_24_port, B => n5850, S => n57, Z
                           => n3376);
   U5168 : MUX2_X1 port map( A => REGISTERS_17_23_port, B => n5851, S => n57, Z
                           => n3375);
   U5169 : MUX2_X1 port map( A => REGISTERS_17_22_port, B => n5852, S => n57, Z
                           => n3374);
   U5170 : MUX2_X1 port map( A => REGISTERS_17_21_port, B => n5853, S => n57, Z
                           => n3373);
   U5171 : MUX2_X1 port map( A => REGISTERS_17_20_port, B => n5854, S => n57, Z
                           => n3372);
   U5172 : MUX2_X1 port map( A => REGISTERS_17_19_port, B => n5855, S => n57, Z
                           => n3371);
   U5173 : MUX2_X1 port map( A => REGISTERS_17_18_port, B => n5856, S => n57, Z
                           => n3370);
   U5174 : MUX2_X1 port map( A => REGISTERS_17_17_port, B => n5857, S => n57, Z
                           => n3369);
   U5175 : MUX2_X1 port map( A => REGISTERS_17_16_port, B => n5858, S => n57, Z
                           => n3368);
   U5176 : MUX2_X1 port map( A => REGISTERS_17_15_port, B => n5859, S => n57, Z
                           => n3367);
   U5177 : MUX2_X1 port map( A => REGISTERS_17_14_port, B => n5860, S => n57, Z
                           => n3366);
   U5178 : MUX2_X1 port map( A => REGISTERS_17_13_port, B => n5861, S => n57, Z
                           => n3365);
   U5179 : MUX2_X1 port map( A => REGISTERS_17_12_port, B => n5862, S => n57, Z
                           => n3364);
   U5180 : MUX2_X1 port map( A => REGISTERS_17_11_port, B => n5863, S => n57, Z
                           => n3363);
   U5181 : MUX2_X1 port map( A => REGISTERS_17_10_port, B => n5864, S => n57, Z
                           => n3362);
   U5182 : MUX2_X1 port map( A => REGISTERS_17_9_port, B => n5865, S => n57, Z 
                           => n3361);
   U5183 : MUX2_X1 port map( A => REGISTERS_17_8_port, B => n5866, S => n57, Z 
                           => n3360);
   U5184 : MUX2_X1 port map( A => REGISTERS_17_7_port, B => n5867, S => n57, Z 
                           => n3359);
   U5185 : MUX2_X1 port map( A => REGISTERS_17_6_port, B => n5868, S => n57, Z 
                           => n3358);
   U5186 : MUX2_X1 port map( A => REGISTERS_17_5_port, B => n5869, S => n57, Z 
                           => n3357);
   U5187 : MUX2_X1 port map( A => REGISTERS_17_4_port, B => n5870, S => n57, Z 
                           => n3356);
   U5188 : MUX2_X1 port map( A => REGISTERS_17_3_port, B => n5871, S => n57, Z 
                           => n3355);
   U5189 : MUX2_X1 port map( A => REGISTERS_17_2_port, B => n5872, S => n57, Z 
                           => n3354);
   U5190 : MUX2_X1 port map( A => REGISTERS_17_1_port, B => n5873, S => n57, Z 
                           => n3353);
   U5191 : MUX2_X1 port map( A => REGISTERS_17_0_port, B => n5874, S => n57, Z 
                           => n3352);
   U5192 : OAI21_X1 port map( B1 => n5878, B2 => n5904, A => n5744, ZN => n5905
                           );
   U5193 : MUX2_X1 port map( A => REGISTERS_18_63_port, B => n5810, S => n59, Z
                           => n3351);
   U5194 : MUX2_X1 port map( A => REGISTERS_18_62_port, B => n5812, S => n59, Z
                           => n3350);
   U5195 : MUX2_X1 port map( A => REGISTERS_18_61_port, B => n5813, S => n59, Z
                           => n3349);
   U5196 : MUX2_X1 port map( A => REGISTERS_18_60_port, B => n5814, S => n59, Z
                           => n3348);
   U5197 : MUX2_X1 port map( A => REGISTERS_18_59_port, B => n5815, S => n59, Z
                           => n3347);
   U5198 : MUX2_X1 port map( A => REGISTERS_18_58_port, B => n5816, S => n59, Z
                           => n3346);
   U5199 : MUX2_X1 port map( A => REGISTERS_18_57_port, B => n5817, S => n59, Z
                           => n3345);
   U5200 : MUX2_X1 port map( A => REGISTERS_18_56_port, B => n5818, S => n59, Z
                           => n3344);
   U5201 : MUX2_X1 port map( A => REGISTERS_18_55_port, B => n5819, S => n59, Z
                           => n3343);
   U5202 : MUX2_X1 port map( A => REGISTERS_18_54_port, B => n5820, S => n59, Z
                           => n3342);
   U5203 : MUX2_X1 port map( A => REGISTERS_18_53_port, B => n5821, S => n59, Z
                           => n3341);
   U5204 : MUX2_X1 port map( A => REGISTERS_18_52_port, B => n5822, S => n59, Z
                           => n3340);
   U5205 : MUX2_X1 port map( A => REGISTERS_18_51_port, B => n5823, S => n59, Z
                           => n3339);
   U5206 : MUX2_X1 port map( A => REGISTERS_18_50_port, B => n5824, S => n59, Z
                           => n3338);
   U5207 : MUX2_X1 port map( A => REGISTERS_18_49_port, B => n5825, S => n59, Z
                           => n3337);
   U5208 : MUX2_X1 port map( A => REGISTERS_18_48_port, B => n5826, S => n59, Z
                           => n3336);
   U5209 : MUX2_X1 port map( A => REGISTERS_18_47_port, B => n5827, S => n59, Z
                           => n3335);
   U5210 : MUX2_X1 port map( A => REGISTERS_18_46_port, B => n5828, S => n59, Z
                           => n3334);
   U5211 : MUX2_X1 port map( A => REGISTERS_18_45_port, B => n5829, S => n59, Z
                           => n3333);
   U5212 : MUX2_X1 port map( A => REGISTERS_18_44_port, B => n5830, S => n59, Z
                           => n3332);
   U5213 : MUX2_X1 port map( A => REGISTERS_18_43_port, B => n5831, S => n59, Z
                           => n3331);
   U5214 : MUX2_X1 port map( A => REGISTERS_18_42_port, B => n5832, S => n59, Z
                           => n3330);
   U5215 : MUX2_X1 port map( A => REGISTERS_18_41_port, B => n5833, S => n59, Z
                           => n3329);
   U5216 : MUX2_X1 port map( A => REGISTERS_18_40_port, B => n5834, S => n59, Z
                           => n3328);
   U5217 : MUX2_X1 port map( A => REGISTERS_18_39_port, B => n5835, S => n59, Z
                           => n3327);
   U5218 : MUX2_X1 port map( A => REGISTERS_18_38_port, B => n5836, S => n59, Z
                           => n3326);
   U5219 : MUX2_X1 port map( A => REGISTERS_18_37_port, B => n5837, S => n59, Z
                           => n3325);
   U5220 : MUX2_X1 port map( A => REGISTERS_18_36_port, B => n5838, S => n59, Z
                           => n3324);
   U5221 : MUX2_X1 port map( A => REGISTERS_18_35_port, B => n5839, S => n59, Z
                           => n3323);
   U5222 : MUX2_X1 port map( A => REGISTERS_18_34_port, B => n5840, S => n59, Z
                           => n3322);
   U5223 : MUX2_X1 port map( A => REGISTERS_18_33_port, B => n5841, S => n59, Z
                           => n3321);
   U5224 : MUX2_X1 port map( A => REGISTERS_18_32_port, B => n5842, S => n59, Z
                           => n3320);
   U5225 : MUX2_X1 port map( A => REGISTERS_18_31_port, B => n5843, S => n59, Z
                           => n3319);
   U5226 : MUX2_X1 port map( A => REGISTERS_18_30_port, B => n5844, S => n59, Z
                           => n3318);
   U5227 : MUX2_X1 port map( A => REGISTERS_18_29_port, B => n5845, S => n59, Z
                           => n3317);
   U5228 : MUX2_X1 port map( A => REGISTERS_18_28_port, B => n5846, S => n59, Z
                           => n3316);
   U5229 : MUX2_X1 port map( A => REGISTERS_18_27_port, B => n5847, S => n59, Z
                           => n3315);
   U5230 : MUX2_X1 port map( A => REGISTERS_18_26_port, B => n5848, S => n59, Z
                           => n3314);
   U5231 : MUX2_X1 port map( A => REGISTERS_18_25_port, B => n5849, S => n59, Z
                           => n3313);
   U5232 : MUX2_X1 port map( A => REGISTERS_18_24_port, B => n5850, S => n59, Z
                           => n3312);
   U5233 : MUX2_X1 port map( A => REGISTERS_18_23_port, B => n5851, S => n59, Z
                           => n3311);
   U5234 : MUX2_X1 port map( A => REGISTERS_18_22_port, B => n5852, S => n59, Z
                           => n3310);
   U5235 : MUX2_X1 port map( A => REGISTERS_18_21_port, B => n5853, S => n59, Z
                           => n3309);
   U5236 : MUX2_X1 port map( A => REGISTERS_18_20_port, B => n5854, S => n59, Z
                           => n3308);
   U5237 : MUX2_X1 port map( A => REGISTERS_18_19_port, B => n5855, S => n59, Z
                           => n3307);
   U5238 : MUX2_X1 port map( A => REGISTERS_18_18_port, B => n5856, S => n59, Z
                           => n3306);
   U5239 : MUX2_X1 port map( A => REGISTERS_18_17_port, B => n5857, S => n59, Z
                           => n3305);
   U5240 : MUX2_X1 port map( A => REGISTERS_18_16_port, B => n5858, S => n59, Z
                           => n3304);
   U5241 : MUX2_X1 port map( A => REGISTERS_18_15_port, B => n5859, S => n59, Z
                           => n3303);
   U5242 : MUX2_X1 port map( A => REGISTERS_18_14_port, B => n5860, S => n59, Z
                           => n3302);
   U5243 : MUX2_X1 port map( A => REGISTERS_18_13_port, B => n5861, S => n59, Z
                           => n3301);
   U5244 : MUX2_X1 port map( A => REGISTERS_18_12_port, B => n5862, S => n59, Z
                           => n3300);
   U5245 : MUX2_X1 port map( A => REGISTERS_18_11_port, B => n5863, S => n59, Z
                           => n3299);
   U5246 : MUX2_X1 port map( A => REGISTERS_18_10_port, B => n5864, S => n59, Z
                           => n3298);
   U5247 : MUX2_X1 port map( A => REGISTERS_18_9_port, B => n5865, S => n59, Z 
                           => n3297);
   U5248 : MUX2_X1 port map( A => REGISTERS_18_8_port, B => n5866, S => n59, Z 
                           => n3296);
   U5249 : MUX2_X1 port map( A => REGISTERS_18_7_port, B => n5867, S => n59, Z 
                           => n3295);
   U5250 : MUX2_X1 port map( A => REGISTERS_18_6_port, B => n5868, S => n59, Z 
                           => n3294);
   U5251 : MUX2_X1 port map( A => REGISTERS_18_5_port, B => n5869, S => n59, Z 
                           => n3293);
   U5252 : MUX2_X1 port map( A => REGISTERS_18_4_port, B => n5870, S => n59, Z 
                           => n3292);
   U5253 : MUX2_X1 port map( A => REGISTERS_18_3_port, B => n5871, S => n59, Z 
                           => n3291);
   U5254 : MUX2_X1 port map( A => REGISTERS_18_2_port, B => n5872, S => n59, Z 
                           => n3290);
   U5255 : MUX2_X1 port map( A => REGISTERS_18_1_port, B => n5873, S => n59, Z 
                           => n3289);
   U5256 : MUX2_X1 port map( A => REGISTERS_18_0_port, B => n5874, S => n59, Z 
                           => n3288);
   U5257 : OAI21_X1 port map( B1 => n5880, B2 => n5904, A => n5744, ZN => n5906
                           );
   U5258 : MUX2_X1 port map( A => REGISTERS_19_63_port, B => n5810, S => n49, Z
                           => n3287);
   U5259 : MUX2_X1 port map( A => REGISTERS_19_62_port, B => n5812, S => n49, Z
                           => n3286);
   U5260 : MUX2_X1 port map( A => REGISTERS_19_61_port, B => n5813, S => n49, Z
                           => n3285);
   U5261 : MUX2_X1 port map( A => REGISTERS_19_60_port, B => n5814, S => n49, Z
                           => n3284);
   U5262 : MUX2_X1 port map( A => REGISTERS_19_59_port, B => n5815, S => n49, Z
                           => n3283);
   U5263 : MUX2_X1 port map( A => REGISTERS_19_58_port, B => n5816, S => n49, Z
                           => n3282);
   U5264 : MUX2_X1 port map( A => REGISTERS_19_57_port, B => n5817, S => n49, Z
                           => n3281);
   U5265 : MUX2_X1 port map( A => REGISTERS_19_56_port, B => n5818, S => n49, Z
                           => n3280);
   U5266 : MUX2_X1 port map( A => REGISTERS_19_55_port, B => n5819, S => n49, Z
                           => n3279);
   U5267 : MUX2_X1 port map( A => REGISTERS_19_54_port, B => n5820, S => n49, Z
                           => n3278);
   U5268 : MUX2_X1 port map( A => REGISTERS_19_53_port, B => n5821, S => n49, Z
                           => n3277);
   U5269 : MUX2_X1 port map( A => REGISTERS_19_52_port, B => n5822, S => n49, Z
                           => n3276);
   U5270 : MUX2_X1 port map( A => REGISTERS_19_51_port, B => n5823, S => n49, Z
                           => n3275);
   U5271 : MUX2_X1 port map( A => REGISTERS_19_50_port, B => n5824, S => n49, Z
                           => n3274);
   U5272 : MUX2_X1 port map( A => REGISTERS_19_49_port, B => n5825, S => n49, Z
                           => n3273);
   U5273 : MUX2_X1 port map( A => REGISTERS_19_48_port, B => n5826, S => n49, Z
                           => n3272);
   U5274 : MUX2_X1 port map( A => REGISTERS_19_47_port, B => n5827, S => n49, Z
                           => n3271);
   U5275 : MUX2_X1 port map( A => REGISTERS_19_46_port, B => n5828, S => n49, Z
                           => n3270);
   U5276 : MUX2_X1 port map( A => REGISTERS_19_45_port, B => n5829, S => n49, Z
                           => n3269);
   U5277 : MUX2_X1 port map( A => REGISTERS_19_44_port, B => n5830, S => n49, Z
                           => n3268);
   U5278 : MUX2_X1 port map( A => REGISTERS_19_43_port, B => n5831, S => n49, Z
                           => n3267);
   U5279 : MUX2_X1 port map( A => REGISTERS_19_42_port, B => n5832, S => n49, Z
                           => n3266);
   U5280 : MUX2_X1 port map( A => REGISTERS_19_41_port, B => n5833, S => n49, Z
                           => n3265);
   U5281 : MUX2_X1 port map( A => REGISTERS_19_40_port, B => n5834, S => n49, Z
                           => n3264);
   U5282 : MUX2_X1 port map( A => REGISTERS_19_39_port, B => n5835, S => n49, Z
                           => n3263);
   U5283 : MUX2_X1 port map( A => REGISTERS_19_38_port, B => n5836, S => n49, Z
                           => n3262);
   U5284 : MUX2_X1 port map( A => REGISTERS_19_37_port, B => n5837, S => n49, Z
                           => n3261);
   U5285 : MUX2_X1 port map( A => REGISTERS_19_36_port, B => n5838, S => n49, Z
                           => n3260);
   U5286 : MUX2_X1 port map( A => REGISTERS_19_35_port, B => n5839, S => n49, Z
                           => n3259);
   U5287 : MUX2_X1 port map( A => REGISTERS_19_34_port, B => n5840, S => n49, Z
                           => n3258);
   U5288 : MUX2_X1 port map( A => REGISTERS_19_33_port, B => n5841, S => n49, Z
                           => n3257);
   U5289 : MUX2_X1 port map( A => REGISTERS_19_32_port, B => n5842, S => n49, Z
                           => n3256);
   U5290 : MUX2_X1 port map( A => REGISTERS_19_31_port, B => n5843, S => n49, Z
                           => n3255);
   U5291 : MUX2_X1 port map( A => REGISTERS_19_30_port, B => n5844, S => n49, Z
                           => n3254);
   U5292 : MUX2_X1 port map( A => REGISTERS_19_29_port, B => n5845, S => n49, Z
                           => n3253);
   U5293 : MUX2_X1 port map( A => REGISTERS_19_28_port, B => n5846, S => n49, Z
                           => n3252);
   U5294 : MUX2_X1 port map( A => REGISTERS_19_27_port, B => n5847, S => n49, Z
                           => n3251);
   U5295 : MUX2_X1 port map( A => REGISTERS_19_26_port, B => n5848, S => n49, Z
                           => n3250);
   U5296 : MUX2_X1 port map( A => REGISTERS_19_25_port, B => n5849, S => n49, Z
                           => n3249);
   U5297 : MUX2_X1 port map( A => REGISTERS_19_24_port, B => n5850, S => n49, Z
                           => n3248);
   U5298 : MUX2_X1 port map( A => REGISTERS_19_23_port, B => n5851, S => n49, Z
                           => n3247);
   U5299 : MUX2_X1 port map( A => REGISTERS_19_22_port, B => n5852, S => n49, Z
                           => n3246);
   U5300 : MUX2_X1 port map( A => REGISTERS_19_21_port, B => n5853, S => n49, Z
                           => n3245);
   U5301 : MUX2_X1 port map( A => REGISTERS_19_20_port, B => n5854, S => n49, Z
                           => n3244);
   U5302 : MUX2_X1 port map( A => REGISTERS_19_19_port, B => n5855, S => n49, Z
                           => n3243);
   U5303 : MUX2_X1 port map( A => REGISTERS_19_18_port, B => n5856, S => n49, Z
                           => n3242);
   U5304 : MUX2_X1 port map( A => REGISTERS_19_17_port, B => n5857, S => n49, Z
                           => n3241);
   U5305 : MUX2_X1 port map( A => REGISTERS_19_16_port, B => n5858, S => n49, Z
                           => n3240);
   U5306 : MUX2_X1 port map( A => REGISTERS_19_15_port, B => n5859, S => n49, Z
                           => n3239);
   U5307 : MUX2_X1 port map( A => REGISTERS_19_14_port, B => n5860, S => n49, Z
                           => n3238);
   U5308 : MUX2_X1 port map( A => REGISTERS_19_13_port, B => n5861, S => n49, Z
                           => n3237);
   U5309 : MUX2_X1 port map( A => REGISTERS_19_12_port, B => n5862, S => n49, Z
                           => n3236);
   U5310 : MUX2_X1 port map( A => REGISTERS_19_11_port, B => n5863, S => n49, Z
                           => n3235);
   U5311 : MUX2_X1 port map( A => REGISTERS_19_10_port, B => n5864, S => n49, Z
                           => n3234);
   U5312 : MUX2_X1 port map( A => REGISTERS_19_9_port, B => n5865, S => n49, Z 
                           => n3233);
   U5313 : MUX2_X1 port map( A => REGISTERS_19_8_port, B => n5866, S => n49, Z 
                           => n3232);
   U5314 : MUX2_X1 port map( A => REGISTERS_19_7_port, B => n5867, S => n49, Z 
                           => n3231);
   U5315 : MUX2_X1 port map( A => REGISTERS_19_6_port, B => n5868, S => n49, Z 
                           => n3230);
   U5316 : MUX2_X1 port map( A => REGISTERS_19_5_port, B => n5869, S => n49, Z 
                           => n3229);
   U5317 : MUX2_X1 port map( A => REGISTERS_19_4_port, B => n5870, S => n49, Z 
                           => n3228);
   U5318 : MUX2_X1 port map( A => REGISTERS_19_3_port, B => n5871, S => n49, Z 
                           => n3227);
   U5319 : MUX2_X1 port map( A => REGISTERS_19_2_port, B => n5872, S => n49, Z 
                           => n3226);
   U5320 : MUX2_X1 port map( A => REGISTERS_19_1_port, B => n5873, S => n49, Z 
                           => n3225);
   U5321 : MUX2_X1 port map( A => REGISTERS_19_0_port, B => n5874, S => n49, Z 
                           => n3224);
   U5322 : OAI21_X1 port map( B1 => n5882, B2 => n5904, A => n5744, ZN => n5907
                           );
   U5323 : MUX2_X1 port map( A => REGISTERS_20_63_port, B => n5810, S => n51, Z
                           => n3223);
   U5324 : MUX2_X1 port map( A => REGISTERS_20_62_port, B => n5812, S => n51, Z
                           => n3222);
   U5325 : MUX2_X1 port map( A => REGISTERS_20_61_port, B => n5813, S => n51, Z
                           => n3221);
   U5326 : MUX2_X1 port map( A => REGISTERS_20_60_port, B => n5814, S => n51, Z
                           => n3220);
   U5327 : MUX2_X1 port map( A => REGISTERS_20_59_port, B => n5815, S => n51, Z
                           => n3219);
   U5328 : MUX2_X1 port map( A => REGISTERS_20_58_port, B => n5816, S => n51, Z
                           => n3218);
   U5329 : MUX2_X1 port map( A => REGISTERS_20_57_port, B => n5817, S => n51, Z
                           => n3217);
   U5330 : MUX2_X1 port map( A => REGISTERS_20_56_port, B => n5818, S => n51, Z
                           => n3216);
   U5331 : MUX2_X1 port map( A => REGISTERS_20_55_port, B => n5819, S => n51, Z
                           => n3215);
   U5332 : MUX2_X1 port map( A => REGISTERS_20_54_port, B => n5820, S => n51, Z
                           => n3214);
   U5333 : MUX2_X1 port map( A => REGISTERS_20_53_port, B => n5821, S => n51, Z
                           => n3213);
   U5334 : MUX2_X1 port map( A => REGISTERS_20_52_port, B => n5822, S => n51, Z
                           => n3212);
   U5335 : MUX2_X1 port map( A => REGISTERS_20_51_port, B => n5823, S => n51, Z
                           => n3211);
   U5336 : MUX2_X1 port map( A => REGISTERS_20_50_port, B => n5824, S => n51, Z
                           => n3210);
   U5337 : MUX2_X1 port map( A => REGISTERS_20_49_port, B => n5825, S => n51, Z
                           => n3209);
   U5338 : MUX2_X1 port map( A => REGISTERS_20_48_port, B => n5826, S => n51, Z
                           => n3208);
   U5339 : MUX2_X1 port map( A => REGISTERS_20_47_port, B => n5827, S => n51, Z
                           => n3207);
   U5340 : MUX2_X1 port map( A => REGISTERS_20_46_port, B => n5828, S => n51, Z
                           => n3206);
   U5341 : MUX2_X1 port map( A => REGISTERS_20_45_port, B => n5829, S => n51, Z
                           => n3205);
   U5342 : MUX2_X1 port map( A => REGISTERS_20_44_port, B => n5830, S => n51, Z
                           => n3204);
   U5343 : MUX2_X1 port map( A => REGISTERS_20_43_port, B => n5831, S => n51, Z
                           => n3203);
   U5344 : MUX2_X1 port map( A => REGISTERS_20_42_port, B => n5832, S => n51, Z
                           => n3202);
   U5345 : MUX2_X1 port map( A => REGISTERS_20_41_port, B => n5833, S => n51, Z
                           => n3201);
   U5346 : MUX2_X1 port map( A => REGISTERS_20_40_port, B => n5834, S => n51, Z
                           => n3200);
   U5347 : MUX2_X1 port map( A => REGISTERS_20_39_port, B => n5835, S => n51, Z
                           => n3199);
   U5348 : MUX2_X1 port map( A => REGISTERS_20_38_port, B => n5836, S => n51, Z
                           => n3198);
   U5349 : MUX2_X1 port map( A => REGISTERS_20_37_port, B => n5837, S => n51, Z
                           => n3197);
   U5350 : MUX2_X1 port map( A => REGISTERS_20_36_port, B => n5838, S => n51, Z
                           => n3196);
   U5351 : MUX2_X1 port map( A => REGISTERS_20_35_port, B => n5839, S => n51, Z
                           => n3195);
   U5352 : MUX2_X1 port map( A => REGISTERS_20_34_port, B => n5840, S => n51, Z
                           => n3194);
   U5353 : MUX2_X1 port map( A => REGISTERS_20_33_port, B => n5841, S => n51, Z
                           => n3193);
   U5354 : MUX2_X1 port map( A => REGISTERS_20_32_port, B => n5842, S => n51, Z
                           => n3192);
   U5355 : MUX2_X1 port map( A => REGISTERS_20_31_port, B => n5843, S => n51, Z
                           => n3191);
   U5356 : MUX2_X1 port map( A => REGISTERS_20_30_port, B => n5844, S => n51, Z
                           => n3190);
   U5357 : MUX2_X1 port map( A => REGISTERS_20_29_port, B => n5845, S => n51, Z
                           => n3189);
   U5358 : MUX2_X1 port map( A => REGISTERS_20_28_port, B => n5846, S => n51, Z
                           => n3188);
   U5359 : MUX2_X1 port map( A => REGISTERS_20_27_port, B => n5847, S => n51, Z
                           => n3187);
   U5360 : MUX2_X1 port map( A => REGISTERS_20_26_port, B => n5848, S => n51, Z
                           => n3186);
   U5361 : MUX2_X1 port map( A => REGISTERS_20_25_port, B => n5849, S => n51, Z
                           => n3185);
   U5362 : MUX2_X1 port map( A => REGISTERS_20_24_port, B => n5850, S => n51, Z
                           => n3184);
   U5363 : MUX2_X1 port map( A => REGISTERS_20_23_port, B => n5851, S => n51, Z
                           => n3183);
   U5364 : MUX2_X1 port map( A => REGISTERS_20_22_port, B => n5852, S => n51, Z
                           => n3182);
   U5365 : MUX2_X1 port map( A => REGISTERS_20_21_port, B => n5853, S => n51, Z
                           => n3181);
   U5366 : MUX2_X1 port map( A => REGISTERS_20_20_port, B => n5854, S => n51, Z
                           => n3180);
   U5367 : MUX2_X1 port map( A => REGISTERS_20_19_port, B => n5855, S => n51, Z
                           => n3179);
   U5368 : MUX2_X1 port map( A => REGISTERS_20_18_port, B => n5856, S => n51, Z
                           => n3178);
   U5369 : MUX2_X1 port map( A => REGISTERS_20_17_port, B => n5857, S => n51, Z
                           => n3177);
   U5370 : MUX2_X1 port map( A => REGISTERS_20_16_port, B => n5858, S => n51, Z
                           => n3176);
   U5371 : MUX2_X1 port map( A => REGISTERS_20_15_port, B => n5859, S => n51, Z
                           => n3175);
   U5372 : MUX2_X1 port map( A => REGISTERS_20_14_port, B => n5860, S => n51, Z
                           => n3174);
   U5373 : MUX2_X1 port map( A => REGISTERS_20_13_port, B => n5861, S => n51, Z
                           => n3173);
   U5374 : MUX2_X1 port map( A => REGISTERS_20_12_port, B => n5862, S => n51, Z
                           => n3172);
   U5375 : MUX2_X1 port map( A => REGISTERS_20_11_port, B => n5863, S => n51, Z
                           => n3171);
   U5376 : MUX2_X1 port map( A => REGISTERS_20_10_port, B => n5864, S => n51, Z
                           => n3170);
   U5377 : MUX2_X1 port map( A => REGISTERS_20_9_port, B => n5865, S => n51, Z 
                           => n3169);
   U5378 : MUX2_X1 port map( A => REGISTERS_20_8_port, B => n5866, S => n51, Z 
                           => n3168);
   U5379 : MUX2_X1 port map( A => REGISTERS_20_7_port, B => n5867, S => n51, Z 
                           => n3167);
   U5380 : MUX2_X1 port map( A => REGISTERS_20_6_port, B => n5868, S => n51, Z 
                           => n3166);
   U5381 : MUX2_X1 port map( A => REGISTERS_20_5_port, B => n5869, S => n51, Z 
                           => n3165);
   U5382 : MUX2_X1 port map( A => REGISTERS_20_4_port, B => n5870, S => n51, Z 
                           => n3164);
   U5383 : MUX2_X1 port map( A => REGISTERS_20_3_port, B => n5871, S => n51, Z 
                           => n3163);
   U5384 : MUX2_X1 port map( A => REGISTERS_20_2_port, B => n5872, S => n51, Z 
                           => n3162);
   U5385 : MUX2_X1 port map( A => REGISTERS_20_1_port, B => n5873, S => n51, Z 
                           => n3161);
   U5386 : MUX2_X1 port map( A => REGISTERS_20_0_port, B => n5874, S => n51, Z 
                           => n3160);
   U5387 : OAI21_X1 port map( B1 => n5884, B2 => n5904, A => n5744, ZN => n5908
                           );
   U5388 : MUX2_X1 port map( A => REGISTERS_21_63_port, B => n5810, S => n45, Z
                           => n3159);
   U5389 : MUX2_X1 port map( A => REGISTERS_21_62_port, B => n5812, S => n45, Z
                           => n3158);
   U5390 : MUX2_X1 port map( A => REGISTERS_21_61_port, B => n5813, S => n45, Z
                           => n3157);
   U5391 : MUX2_X1 port map( A => REGISTERS_21_60_port, B => n5814, S => n45, Z
                           => n3156);
   U5392 : MUX2_X1 port map( A => REGISTERS_21_59_port, B => n5815, S => n45, Z
                           => n3155);
   U5393 : MUX2_X1 port map( A => REGISTERS_21_58_port, B => n5816, S => n45, Z
                           => n3154);
   U5394 : MUX2_X1 port map( A => REGISTERS_21_57_port, B => n5817, S => n45, Z
                           => n3153);
   U5395 : MUX2_X1 port map( A => REGISTERS_21_56_port, B => n5818, S => n45, Z
                           => n3152);
   U5396 : MUX2_X1 port map( A => REGISTERS_21_55_port, B => n5819, S => n45, Z
                           => n3151);
   U5397 : MUX2_X1 port map( A => REGISTERS_21_54_port, B => n5820, S => n45, Z
                           => n3150);
   U5398 : MUX2_X1 port map( A => REGISTERS_21_53_port, B => n5821, S => n45, Z
                           => n3149);
   U5399 : MUX2_X1 port map( A => REGISTERS_21_52_port, B => n5822, S => n45, Z
                           => n3148);
   U5400 : MUX2_X1 port map( A => REGISTERS_21_51_port, B => n5823, S => n45, Z
                           => n3147);
   U5401 : MUX2_X1 port map( A => REGISTERS_21_50_port, B => n5824, S => n45, Z
                           => n3146);
   U5402 : MUX2_X1 port map( A => REGISTERS_21_49_port, B => n5825, S => n45, Z
                           => n3145);
   U5403 : MUX2_X1 port map( A => REGISTERS_21_48_port, B => n5826, S => n45, Z
                           => n3144);
   U5404 : MUX2_X1 port map( A => REGISTERS_21_47_port, B => n5827, S => n45, Z
                           => n3143);
   U5405 : MUX2_X1 port map( A => REGISTERS_21_46_port, B => n5828, S => n45, Z
                           => n3142);
   U5406 : MUX2_X1 port map( A => REGISTERS_21_45_port, B => n5829, S => n45, Z
                           => n3141);
   U5407 : MUX2_X1 port map( A => REGISTERS_21_44_port, B => n5830, S => n45, Z
                           => n3140);
   U5408 : MUX2_X1 port map( A => REGISTERS_21_43_port, B => n5831, S => n45, Z
                           => n3139);
   U5409 : MUX2_X1 port map( A => REGISTERS_21_42_port, B => n5832, S => n45, Z
                           => n3138);
   U5410 : MUX2_X1 port map( A => REGISTERS_21_41_port, B => n5833, S => n45, Z
                           => n3137);
   U5411 : MUX2_X1 port map( A => REGISTERS_21_40_port, B => n5834, S => n45, Z
                           => n3136);
   U5412 : MUX2_X1 port map( A => REGISTERS_21_39_port, B => n5835, S => n45, Z
                           => n3135);
   U5413 : MUX2_X1 port map( A => REGISTERS_21_38_port, B => n5836, S => n45, Z
                           => n3134);
   U5414 : MUX2_X1 port map( A => REGISTERS_21_37_port, B => n5837, S => n45, Z
                           => n3133);
   U5415 : MUX2_X1 port map( A => REGISTERS_21_36_port, B => n5838, S => n45, Z
                           => n3132);
   U5416 : MUX2_X1 port map( A => REGISTERS_21_35_port, B => n5839, S => n45, Z
                           => n3131);
   U5417 : MUX2_X1 port map( A => REGISTERS_21_34_port, B => n5840, S => n45, Z
                           => n3130);
   U5418 : MUX2_X1 port map( A => REGISTERS_21_33_port, B => n5841, S => n45, Z
                           => n3129);
   U5419 : MUX2_X1 port map( A => REGISTERS_21_32_port, B => n5842, S => n45, Z
                           => n3128);
   U5420 : MUX2_X1 port map( A => REGISTERS_21_31_port, B => n5843, S => n45, Z
                           => n3127);
   U5421 : MUX2_X1 port map( A => REGISTERS_21_30_port, B => n5844, S => n45, Z
                           => n3126);
   U5422 : MUX2_X1 port map( A => REGISTERS_21_29_port, B => n5845, S => n45, Z
                           => n3125);
   U5423 : MUX2_X1 port map( A => REGISTERS_21_28_port, B => n5846, S => n45, Z
                           => n3124);
   U5424 : MUX2_X1 port map( A => REGISTERS_21_27_port, B => n5847, S => n45, Z
                           => n3123);
   U5425 : MUX2_X1 port map( A => REGISTERS_21_26_port, B => n5848, S => n45, Z
                           => n3122);
   U5426 : MUX2_X1 port map( A => REGISTERS_21_25_port, B => n5849, S => n45, Z
                           => n3121);
   U5427 : MUX2_X1 port map( A => REGISTERS_21_24_port, B => n5850, S => n45, Z
                           => n3120);
   U5428 : MUX2_X1 port map( A => REGISTERS_21_23_port, B => n5851, S => n45, Z
                           => n3119);
   U5429 : MUX2_X1 port map( A => REGISTERS_21_22_port, B => n5852, S => n45, Z
                           => n3118);
   U5430 : MUX2_X1 port map( A => REGISTERS_21_21_port, B => n5853, S => n45, Z
                           => n3117);
   U5431 : MUX2_X1 port map( A => REGISTERS_21_20_port, B => n5854, S => n45, Z
                           => n3116);
   U5432 : MUX2_X1 port map( A => REGISTERS_21_19_port, B => n5855, S => n45, Z
                           => n3115);
   U5433 : MUX2_X1 port map( A => REGISTERS_21_18_port, B => n5856, S => n45, Z
                           => n3114);
   U5434 : MUX2_X1 port map( A => REGISTERS_21_17_port, B => n5857, S => n45, Z
                           => n3113);
   U5435 : MUX2_X1 port map( A => REGISTERS_21_16_port, B => n5858, S => n45, Z
                           => n3112);
   U5436 : MUX2_X1 port map( A => REGISTERS_21_15_port, B => n5859, S => n45, Z
                           => n3111);
   U5437 : MUX2_X1 port map( A => REGISTERS_21_14_port, B => n5860, S => n45, Z
                           => n3110);
   U5438 : MUX2_X1 port map( A => REGISTERS_21_13_port, B => n5861, S => n45, Z
                           => n3109);
   U5439 : MUX2_X1 port map( A => REGISTERS_21_12_port, B => n5862, S => n45, Z
                           => n3108);
   U5440 : MUX2_X1 port map( A => REGISTERS_21_11_port, B => n5863, S => n45, Z
                           => n3107);
   U5441 : MUX2_X1 port map( A => REGISTERS_21_10_port, B => n5864, S => n45, Z
                           => n3106);
   U5442 : MUX2_X1 port map( A => REGISTERS_21_9_port, B => n5865, S => n45, Z 
                           => n3105);
   U5443 : MUX2_X1 port map( A => REGISTERS_21_8_port, B => n5866, S => n45, Z 
                           => n3104);
   U5444 : MUX2_X1 port map( A => REGISTERS_21_7_port, B => n5867, S => n45, Z 
                           => n3103);
   U5445 : MUX2_X1 port map( A => REGISTERS_21_6_port, B => n5868, S => n45, Z 
                           => n3102);
   U5446 : MUX2_X1 port map( A => REGISTERS_21_5_port, B => n5869, S => n45, Z 
                           => n3101);
   U5447 : MUX2_X1 port map( A => REGISTERS_21_4_port, B => n5870, S => n45, Z 
                           => n3100);
   U5448 : MUX2_X1 port map( A => REGISTERS_21_3_port, B => n5871, S => n45, Z 
                           => n3099);
   U5449 : MUX2_X1 port map( A => REGISTERS_21_2_port, B => n5872, S => n45, Z 
                           => n3098);
   U5450 : MUX2_X1 port map( A => REGISTERS_21_1_port, B => n5873, S => n45, Z 
                           => n3097);
   U5451 : MUX2_X1 port map( A => REGISTERS_21_0_port, B => n5874, S => n45, Z 
                           => n3096);
   U5452 : OAI21_X1 port map( B1 => n5886, B2 => n5904, A => n5744, ZN => n5909
                           );
   U5453 : MUX2_X1 port map( A => REGISTERS_22_63_port, B => n5810, S => n47, Z
                           => n3095);
   U5454 : MUX2_X1 port map( A => REGISTERS_22_62_port, B => n5812, S => n47, Z
                           => n3094);
   U5455 : MUX2_X1 port map( A => REGISTERS_22_61_port, B => n5813, S => n47, Z
                           => n3093);
   U5456 : MUX2_X1 port map( A => REGISTERS_22_60_port, B => n5814, S => n47, Z
                           => n3092);
   U5457 : MUX2_X1 port map( A => REGISTERS_22_59_port, B => n5815, S => n47, Z
                           => n3091);
   U5458 : MUX2_X1 port map( A => REGISTERS_22_58_port, B => n5816, S => n47, Z
                           => n3090);
   U5459 : MUX2_X1 port map( A => REGISTERS_22_57_port, B => n5817, S => n47, Z
                           => n3089);
   U5460 : MUX2_X1 port map( A => REGISTERS_22_56_port, B => n5818, S => n47, Z
                           => n3088);
   U5461 : MUX2_X1 port map( A => REGISTERS_22_55_port, B => n5819, S => n47, Z
                           => n3087);
   U5462 : MUX2_X1 port map( A => REGISTERS_22_54_port, B => n5820, S => n47, Z
                           => n3086);
   U5463 : MUX2_X1 port map( A => REGISTERS_22_53_port, B => n5821, S => n47, Z
                           => n3085);
   U5464 : MUX2_X1 port map( A => REGISTERS_22_52_port, B => n5822, S => n47, Z
                           => n3084);
   U5465 : MUX2_X1 port map( A => REGISTERS_22_51_port, B => n5823, S => n47, Z
                           => n3083);
   U5466 : MUX2_X1 port map( A => REGISTERS_22_50_port, B => n5824, S => n47, Z
                           => n3082);
   U5467 : MUX2_X1 port map( A => REGISTERS_22_49_port, B => n5825, S => n47, Z
                           => n3081);
   U5468 : MUX2_X1 port map( A => REGISTERS_22_48_port, B => n5826, S => n47, Z
                           => n3080);
   U5469 : MUX2_X1 port map( A => REGISTERS_22_47_port, B => n5827, S => n47, Z
                           => n3079);
   U5470 : MUX2_X1 port map( A => REGISTERS_22_46_port, B => n5828, S => n47, Z
                           => n3078);
   U5471 : MUX2_X1 port map( A => REGISTERS_22_45_port, B => n5829, S => n47, Z
                           => n3077);
   U5472 : MUX2_X1 port map( A => REGISTERS_22_44_port, B => n5830, S => n47, Z
                           => n3076);
   U5473 : MUX2_X1 port map( A => REGISTERS_22_43_port, B => n5831, S => n47, Z
                           => n3075);
   U5474 : MUX2_X1 port map( A => REGISTERS_22_42_port, B => n5832, S => n47, Z
                           => n3074);
   U5475 : MUX2_X1 port map( A => REGISTERS_22_41_port, B => n5833, S => n47, Z
                           => n3073);
   U5476 : MUX2_X1 port map( A => REGISTERS_22_40_port, B => n5834, S => n47, Z
                           => n3072);
   U5477 : MUX2_X1 port map( A => REGISTERS_22_39_port, B => n5835, S => n47, Z
                           => n3071);
   U5478 : MUX2_X1 port map( A => REGISTERS_22_38_port, B => n5836, S => n47, Z
                           => n3070);
   U5479 : MUX2_X1 port map( A => REGISTERS_22_37_port, B => n5837, S => n47, Z
                           => n3069);
   U5480 : MUX2_X1 port map( A => REGISTERS_22_36_port, B => n5838, S => n47, Z
                           => n3068);
   U5481 : MUX2_X1 port map( A => REGISTERS_22_35_port, B => n5839, S => n47, Z
                           => n3067);
   U5482 : MUX2_X1 port map( A => REGISTERS_22_34_port, B => n5840, S => n47, Z
                           => n3066);
   U5483 : MUX2_X1 port map( A => REGISTERS_22_33_port, B => n5841, S => n47, Z
                           => n3065);
   U5484 : MUX2_X1 port map( A => REGISTERS_22_32_port, B => n5842, S => n47, Z
                           => n3064);
   U5485 : MUX2_X1 port map( A => REGISTERS_22_31_port, B => n5843, S => n47, Z
                           => n3063);
   U5486 : MUX2_X1 port map( A => REGISTERS_22_30_port, B => n5844, S => n47, Z
                           => n3062);
   U5487 : MUX2_X1 port map( A => REGISTERS_22_29_port, B => n5845, S => n47, Z
                           => n3061);
   U5488 : MUX2_X1 port map( A => REGISTERS_22_28_port, B => n5846, S => n47, Z
                           => n3060);
   U5489 : MUX2_X1 port map( A => REGISTERS_22_27_port, B => n5847, S => n47, Z
                           => n3059);
   U5490 : MUX2_X1 port map( A => REGISTERS_22_26_port, B => n5848, S => n47, Z
                           => n3058);
   U5491 : MUX2_X1 port map( A => REGISTERS_22_25_port, B => n5849, S => n47, Z
                           => n3057);
   U5492 : MUX2_X1 port map( A => REGISTERS_22_24_port, B => n5850, S => n47, Z
                           => n3056);
   U5493 : MUX2_X1 port map( A => REGISTERS_22_23_port, B => n5851, S => n47, Z
                           => n3055);
   U5494 : MUX2_X1 port map( A => REGISTERS_22_22_port, B => n5852, S => n47, Z
                           => n3054);
   U5495 : MUX2_X1 port map( A => REGISTERS_22_21_port, B => n5853, S => n47, Z
                           => n3053);
   U5496 : MUX2_X1 port map( A => REGISTERS_22_20_port, B => n5854, S => n47, Z
                           => n3052);
   U5497 : MUX2_X1 port map( A => REGISTERS_22_19_port, B => n5855, S => n47, Z
                           => n3051);
   U5498 : MUX2_X1 port map( A => REGISTERS_22_18_port, B => n5856, S => n47, Z
                           => n3050);
   U5499 : MUX2_X1 port map( A => REGISTERS_22_17_port, B => n5857, S => n47, Z
                           => n3049);
   U5500 : MUX2_X1 port map( A => REGISTERS_22_16_port, B => n5858, S => n47, Z
                           => n3048);
   U5501 : MUX2_X1 port map( A => REGISTERS_22_15_port, B => n5859, S => n47, Z
                           => n3047);
   U5502 : MUX2_X1 port map( A => REGISTERS_22_14_port, B => n5860, S => n47, Z
                           => n3046);
   U5503 : MUX2_X1 port map( A => REGISTERS_22_13_port, B => n5861, S => n47, Z
                           => n3045);
   U5504 : MUX2_X1 port map( A => REGISTERS_22_12_port, B => n5862, S => n47, Z
                           => n3044);
   U5505 : MUX2_X1 port map( A => REGISTERS_22_11_port, B => n5863, S => n47, Z
                           => n3043);
   U5506 : MUX2_X1 port map( A => REGISTERS_22_10_port, B => n5864, S => n47, Z
                           => n3042);
   U5507 : MUX2_X1 port map( A => REGISTERS_22_9_port, B => n5865, S => n47, Z 
                           => n3041);
   U5508 : MUX2_X1 port map( A => REGISTERS_22_8_port, B => n5866, S => n47, Z 
                           => n3040);
   U5509 : MUX2_X1 port map( A => REGISTERS_22_7_port, B => n5867, S => n47, Z 
                           => n3039);
   U5510 : MUX2_X1 port map( A => REGISTERS_22_6_port, B => n5868, S => n47, Z 
                           => n3038);
   U5511 : MUX2_X1 port map( A => REGISTERS_22_5_port, B => n5869, S => n47, Z 
                           => n3037);
   U5512 : MUX2_X1 port map( A => REGISTERS_22_4_port, B => n5870, S => n47, Z 
                           => n3036);
   U5513 : MUX2_X1 port map( A => REGISTERS_22_3_port, B => n5871, S => n47, Z 
                           => n3035);
   U5514 : MUX2_X1 port map( A => REGISTERS_22_2_port, B => n5872, S => n47, Z 
                           => n3034);
   U5515 : MUX2_X1 port map( A => REGISTERS_22_1_port, B => n5873, S => n47, Z 
                           => n3033);
   U5516 : MUX2_X1 port map( A => REGISTERS_22_0_port, B => n5874, S => n47, Z 
                           => n3032);
   U5517 : OAI21_X1 port map( B1 => n5888, B2 => n5904, A => n5744, ZN => n5910
                           );
   U5518 : MUX2_X1 port map( A => REGISTERS_23_63_port, B => n5810, S => n41, Z
                           => n3031);
   U5519 : MUX2_X1 port map( A => REGISTERS_23_62_port, B => n5812, S => n41, Z
                           => n3030);
   U5520 : MUX2_X1 port map( A => REGISTERS_23_61_port, B => n5813, S => n41, Z
                           => n3029);
   U5521 : MUX2_X1 port map( A => REGISTERS_23_60_port, B => n5814, S => n41, Z
                           => n3028);
   U5522 : MUX2_X1 port map( A => REGISTERS_23_59_port, B => n5815, S => n41, Z
                           => n3027);
   U5523 : MUX2_X1 port map( A => REGISTERS_23_58_port, B => n5816, S => n41, Z
                           => n3026);
   U5524 : MUX2_X1 port map( A => REGISTERS_23_57_port, B => n5817, S => n41, Z
                           => n3025);
   U5525 : MUX2_X1 port map( A => REGISTERS_23_56_port, B => n5818, S => n41, Z
                           => n3024);
   U5526 : MUX2_X1 port map( A => REGISTERS_23_55_port, B => n5819, S => n41, Z
                           => n3023);
   U5527 : MUX2_X1 port map( A => REGISTERS_23_54_port, B => n5820, S => n41, Z
                           => n3022);
   U5528 : MUX2_X1 port map( A => REGISTERS_23_53_port, B => n5821, S => n41, Z
                           => n3021);
   U5529 : MUX2_X1 port map( A => REGISTERS_23_52_port, B => n5822, S => n41, Z
                           => n3020);
   U5530 : MUX2_X1 port map( A => REGISTERS_23_51_port, B => n5823, S => n41, Z
                           => n3019);
   U5531 : MUX2_X1 port map( A => REGISTERS_23_50_port, B => n5824, S => n41, Z
                           => n3018);
   U5532 : MUX2_X1 port map( A => REGISTERS_23_49_port, B => n5825, S => n41, Z
                           => n3017);
   U5533 : MUX2_X1 port map( A => REGISTERS_23_48_port, B => n5826, S => n41, Z
                           => n3016);
   U5534 : MUX2_X1 port map( A => REGISTERS_23_47_port, B => n5827, S => n41, Z
                           => n3015);
   U5535 : MUX2_X1 port map( A => REGISTERS_23_46_port, B => n5828, S => n41, Z
                           => n3014);
   U5536 : MUX2_X1 port map( A => REGISTERS_23_45_port, B => n5829, S => n41, Z
                           => n3013);
   U5537 : MUX2_X1 port map( A => REGISTERS_23_44_port, B => n5830, S => n41, Z
                           => n3012);
   U5538 : MUX2_X1 port map( A => REGISTERS_23_43_port, B => n5831, S => n41, Z
                           => n3011);
   U5539 : MUX2_X1 port map( A => REGISTERS_23_42_port, B => n5832, S => n41, Z
                           => n3010);
   U5540 : MUX2_X1 port map( A => REGISTERS_23_41_port, B => n5833, S => n41, Z
                           => n3009);
   U5541 : MUX2_X1 port map( A => REGISTERS_23_40_port, B => n5834, S => n41, Z
                           => n3008);
   U5542 : MUX2_X1 port map( A => REGISTERS_23_39_port, B => n5835, S => n41, Z
                           => n3007);
   U5543 : MUX2_X1 port map( A => REGISTERS_23_38_port, B => n5836, S => n41, Z
                           => n3006);
   U5544 : MUX2_X1 port map( A => REGISTERS_23_37_port, B => n5837, S => n41, Z
                           => n3005);
   U5545 : MUX2_X1 port map( A => REGISTERS_23_36_port, B => n5838, S => n41, Z
                           => n3004);
   U5546 : MUX2_X1 port map( A => REGISTERS_23_35_port, B => n5839, S => n41, Z
                           => n3003);
   U5547 : MUX2_X1 port map( A => REGISTERS_23_34_port, B => n5840, S => n41, Z
                           => n3002);
   U5548 : MUX2_X1 port map( A => REGISTERS_23_33_port, B => n5841, S => n41, Z
                           => n3001);
   U5549 : MUX2_X1 port map( A => REGISTERS_23_32_port, B => n5842, S => n41, Z
                           => n3000);
   U5550 : MUX2_X1 port map( A => REGISTERS_23_31_port, B => n5843, S => n41, Z
                           => n2999);
   U5551 : MUX2_X1 port map( A => REGISTERS_23_30_port, B => n5844, S => n41, Z
                           => n2998);
   U5552 : MUX2_X1 port map( A => REGISTERS_23_29_port, B => n5845, S => n41, Z
                           => n2997);
   U5553 : MUX2_X1 port map( A => REGISTERS_23_28_port, B => n5846, S => n41, Z
                           => n2996);
   U5554 : MUX2_X1 port map( A => REGISTERS_23_27_port, B => n5847, S => n41, Z
                           => n2995);
   U5555 : MUX2_X1 port map( A => REGISTERS_23_26_port, B => n5848, S => n41, Z
                           => n2994);
   U5556 : MUX2_X1 port map( A => REGISTERS_23_25_port, B => n5849, S => n41, Z
                           => n2993);
   U5557 : MUX2_X1 port map( A => REGISTERS_23_24_port, B => n5850, S => n41, Z
                           => n2992);
   U5558 : MUX2_X1 port map( A => REGISTERS_23_23_port, B => n5851, S => n41, Z
                           => n2991);
   U5559 : MUX2_X1 port map( A => REGISTERS_23_22_port, B => n5852, S => n41, Z
                           => n2990);
   U5560 : MUX2_X1 port map( A => REGISTERS_23_21_port, B => n5853, S => n41, Z
                           => n2989);
   U5561 : MUX2_X1 port map( A => REGISTERS_23_20_port, B => n5854, S => n41, Z
                           => n2988);
   U5562 : MUX2_X1 port map( A => REGISTERS_23_19_port, B => n5855, S => n41, Z
                           => n2987);
   U5563 : MUX2_X1 port map( A => REGISTERS_23_18_port, B => n5856, S => n41, Z
                           => n2986);
   U5564 : MUX2_X1 port map( A => REGISTERS_23_17_port, B => n5857, S => n41, Z
                           => n2985);
   U5565 : MUX2_X1 port map( A => REGISTERS_23_16_port, B => n5858, S => n41, Z
                           => n2984);
   U5566 : MUX2_X1 port map( A => REGISTERS_23_15_port, B => n5859, S => n41, Z
                           => n2983);
   U5567 : MUX2_X1 port map( A => REGISTERS_23_14_port, B => n5860, S => n41, Z
                           => n2982);
   U5568 : MUX2_X1 port map( A => REGISTERS_23_13_port, B => n5861, S => n41, Z
                           => n2981);
   U5569 : MUX2_X1 port map( A => REGISTERS_23_12_port, B => n5862, S => n41, Z
                           => n2980);
   U5570 : MUX2_X1 port map( A => REGISTERS_23_11_port, B => n5863, S => n41, Z
                           => n2979);
   U5571 : MUX2_X1 port map( A => REGISTERS_23_10_port, B => n5864, S => n41, Z
                           => n2978);
   U5572 : MUX2_X1 port map( A => REGISTERS_23_9_port, B => n5865, S => n41, Z 
                           => n2977);
   U5573 : MUX2_X1 port map( A => REGISTERS_23_8_port, B => n5866, S => n41, Z 
                           => n2976);
   U5574 : MUX2_X1 port map( A => REGISTERS_23_7_port, B => n5867, S => n41, Z 
                           => n2975);
   U5575 : MUX2_X1 port map( A => REGISTERS_23_6_port, B => n5868, S => n41, Z 
                           => n2974);
   U5576 : MUX2_X1 port map( A => REGISTERS_23_5_port, B => n5869, S => n41, Z 
                           => n2973);
   U5577 : MUX2_X1 port map( A => REGISTERS_23_4_port, B => n5870, S => n41, Z 
                           => n2972);
   U5578 : MUX2_X1 port map( A => REGISTERS_23_3_port, B => n5871, S => n41, Z 
                           => n2971);
   U5579 : MUX2_X1 port map( A => REGISTERS_23_2_port, B => n5872, S => n41, Z 
                           => n2970);
   U5580 : MUX2_X1 port map( A => REGISTERS_23_1_port, B => n5873, S => n41, Z 
                           => n2969);
   U5581 : MUX2_X1 port map( A => REGISTERS_23_0_port, B => n5874, S => n41, Z 
                           => n2968);
   U5582 : OAI21_X1 port map( B1 => n5890, B2 => n5904, A => n5744, ZN => n5911
                           );
   U5583 : NAND3_X1 port map( A1 => n5893, A2 => n5891, A3 => ADD_WR(4), ZN => 
                           n5904);
   U5584 : INV_X1 port map( A => ADD_WR(3), ZN => n5891);
   U5585 : MUX2_X1 port map( A => REGISTERS_24_63_port, B => n5810, S => n43, Z
                           => n2967);
   U5586 : MUX2_X1 port map( A => REGISTERS_24_62_port, B => n5812, S => n43, Z
                           => n2966);
   U5587 : MUX2_X1 port map( A => REGISTERS_24_61_port, B => n5813, S => n43, Z
                           => n2965);
   U5588 : MUX2_X1 port map( A => REGISTERS_24_60_port, B => n5814, S => n43, Z
                           => n2964);
   U5589 : MUX2_X1 port map( A => REGISTERS_24_59_port, B => n5815, S => n43, Z
                           => n2963);
   U5590 : MUX2_X1 port map( A => REGISTERS_24_58_port, B => n5816, S => n43, Z
                           => n2962);
   U5591 : MUX2_X1 port map( A => REGISTERS_24_57_port, B => n5817, S => n43, Z
                           => n2961);
   U5592 : MUX2_X1 port map( A => REGISTERS_24_56_port, B => n5818, S => n43, Z
                           => n2960);
   U5593 : MUX2_X1 port map( A => REGISTERS_24_55_port, B => n5819, S => n43, Z
                           => n2959);
   U5594 : MUX2_X1 port map( A => REGISTERS_24_54_port, B => n5820, S => n43, Z
                           => n2958);
   U5595 : MUX2_X1 port map( A => REGISTERS_24_53_port, B => n5821, S => n43, Z
                           => n2957);
   U5596 : MUX2_X1 port map( A => REGISTERS_24_52_port, B => n5822, S => n43, Z
                           => n2956);
   U5597 : MUX2_X1 port map( A => REGISTERS_24_51_port, B => n5823, S => n43, Z
                           => n2955);
   U5598 : MUX2_X1 port map( A => REGISTERS_24_50_port, B => n5824, S => n43, Z
                           => n2954);
   U5599 : MUX2_X1 port map( A => REGISTERS_24_49_port, B => n5825, S => n43, Z
                           => n2953);
   U5600 : MUX2_X1 port map( A => REGISTERS_24_48_port, B => n5826, S => n43, Z
                           => n2952);
   U5601 : MUX2_X1 port map( A => REGISTERS_24_47_port, B => n5827, S => n43, Z
                           => n2951);
   U5602 : MUX2_X1 port map( A => REGISTERS_24_46_port, B => n5828, S => n43, Z
                           => n2950);
   U5603 : MUX2_X1 port map( A => REGISTERS_24_45_port, B => n5829, S => n43, Z
                           => n2949);
   U5604 : MUX2_X1 port map( A => REGISTERS_24_44_port, B => n5830, S => n43, Z
                           => n2948);
   U5605 : MUX2_X1 port map( A => REGISTERS_24_43_port, B => n5831, S => n43, Z
                           => n2947);
   U5606 : MUX2_X1 port map( A => REGISTERS_24_42_port, B => n5832, S => n43, Z
                           => n2946);
   U5607 : MUX2_X1 port map( A => REGISTERS_24_41_port, B => n5833, S => n43, Z
                           => n2945);
   U5608 : MUX2_X1 port map( A => REGISTERS_24_40_port, B => n5834, S => n43, Z
                           => n2944);
   U5609 : MUX2_X1 port map( A => REGISTERS_24_39_port, B => n5835, S => n43, Z
                           => n2943);
   U5610 : MUX2_X1 port map( A => REGISTERS_24_38_port, B => n5836, S => n43, Z
                           => n2942);
   U5611 : MUX2_X1 port map( A => REGISTERS_24_37_port, B => n5837, S => n43, Z
                           => n2941);
   U5612 : MUX2_X1 port map( A => REGISTERS_24_36_port, B => n5838, S => n43, Z
                           => n2940);
   U5613 : MUX2_X1 port map( A => REGISTERS_24_35_port, B => n5839, S => n43, Z
                           => n2939);
   U5614 : MUX2_X1 port map( A => REGISTERS_24_34_port, B => n5840, S => n43, Z
                           => n2938);
   U5615 : MUX2_X1 port map( A => REGISTERS_24_33_port, B => n5841, S => n43, Z
                           => n2937);
   U5616 : MUX2_X1 port map( A => REGISTERS_24_32_port, B => n5842, S => n43, Z
                           => n2936);
   U5617 : MUX2_X1 port map( A => REGISTERS_24_31_port, B => n5843, S => n43, Z
                           => n2935);
   U5618 : MUX2_X1 port map( A => REGISTERS_24_30_port, B => n5844, S => n43, Z
                           => n2934);
   U5619 : MUX2_X1 port map( A => REGISTERS_24_29_port, B => n5845, S => n43, Z
                           => n2933);
   U5620 : MUX2_X1 port map( A => REGISTERS_24_28_port, B => n5846, S => n43, Z
                           => n2932);
   U5621 : MUX2_X1 port map( A => REGISTERS_24_27_port, B => n5847, S => n43, Z
                           => n2931);
   U5622 : MUX2_X1 port map( A => REGISTERS_24_26_port, B => n5848, S => n43, Z
                           => n2930);
   U5623 : MUX2_X1 port map( A => REGISTERS_24_25_port, B => n5849, S => n43, Z
                           => n2929);
   U5624 : MUX2_X1 port map( A => REGISTERS_24_24_port, B => n5850, S => n43, Z
                           => n2928);
   U5625 : MUX2_X1 port map( A => REGISTERS_24_23_port, B => n5851, S => n43, Z
                           => n2927);
   U5626 : MUX2_X1 port map( A => REGISTERS_24_22_port, B => n5852, S => n43, Z
                           => n2926);
   U5627 : MUX2_X1 port map( A => REGISTERS_24_21_port, B => n5853, S => n43, Z
                           => n2925);
   U5628 : MUX2_X1 port map( A => REGISTERS_24_20_port, B => n5854, S => n43, Z
                           => n2924);
   U5629 : MUX2_X1 port map( A => REGISTERS_24_19_port, B => n5855, S => n43, Z
                           => n2923);
   U5630 : MUX2_X1 port map( A => REGISTERS_24_18_port, B => n5856, S => n43, Z
                           => n2922);
   U5631 : MUX2_X1 port map( A => REGISTERS_24_17_port, B => n5857, S => n43, Z
                           => n2921);
   U5632 : MUX2_X1 port map( A => REGISTERS_24_16_port, B => n5858, S => n43, Z
                           => n2920);
   U5633 : MUX2_X1 port map( A => REGISTERS_24_15_port, B => n5859, S => n43, Z
                           => n2919);
   U5634 : MUX2_X1 port map( A => REGISTERS_24_14_port, B => n5860, S => n43, Z
                           => n2918);
   U5635 : MUX2_X1 port map( A => REGISTERS_24_13_port, B => n5861, S => n43, Z
                           => n2917);
   U5636 : MUX2_X1 port map( A => REGISTERS_24_12_port, B => n5862, S => n43, Z
                           => n2916);
   U5637 : MUX2_X1 port map( A => REGISTERS_24_11_port, B => n5863, S => n43, Z
                           => n2915);
   U5638 : MUX2_X1 port map( A => REGISTERS_24_10_port, B => n5864, S => n43, Z
                           => n2914);
   U5639 : MUX2_X1 port map( A => REGISTERS_24_9_port, B => n5865, S => n43, Z 
                           => n2913);
   U5640 : MUX2_X1 port map( A => REGISTERS_24_8_port, B => n5866, S => n43, Z 
                           => n2912);
   U5641 : MUX2_X1 port map( A => REGISTERS_24_7_port, B => n5867, S => n43, Z 
                           => n2911);
   U5642 : MUX2_X1 port map( A => REGISTERS_24_6_port, B => n5868, S => n43, Z 
                           => n2910);
   U5643 : MUX2_X1 port map( A => REGISTERS_24_5_port, B => n5869, S => n43, Z 
                           => n2909);
   U5644 : MUX2_X1 port map( A => REGISTERS_24_4_port, B => n5870, S => n43, Z 
                           => n2908);
   U5645 : MUX2_X1 port map( A => REGISTERS_24_3_port, B => n5871, S => n43, Z 
                           => n2907);
   U5646 : MUX2_X1 port map( A => REGISTERS_24_2_port, B => n5872, S => n43, Z 
                           => n2906);
   U5647 : MUX2_X1 port map( A => REGISTERS_24_1_port, B => n5873, S => n43, Z 
                           => n2905);
   U5648 : MUX2_X1 port map( A => REGISTERS_24_0_port, B => n5874, S => n43, Z 
                           => n2904);
   U5649 : OAI21_X1 port map( B1 => n5876, B2 => n5913, A => n5744, ZN => n5912
                           );
   U5650 : NAND3_X1 port map( A1 => n5914, A2 => n5915, A3 => n5916, ZN => 
                           n5876);
   U5651 : MUX2_X1 port map( A => REGISTERS_25_63_port, B => n5810, S => n37, Z
                           => n2903);
   U5652 : MUX2_X1 port map( A => REGISTERS_25_62_port, B => n5812, S => n37, Z
                           => n2902);
   U5653 : MUX2_X1 port map( A => REGISTERS_25_61_port, B => n5813, S => n37, Z
                           => n2901);
   U5654 : MUX2_X1 port map( A => REGISTERS_25_60_port, B => n5814, S => n37, Z
                           => n2900);
   U5655 : MUX2_X1 port map( A => REGISTERS_25_59_port, B => n5815, S => n37, Z
                           => n2899);
   U5656 : MUX2_X1 port map( A => REGISTERS_25_58_port, B => n5816, S => n37, Z
                           => n2898);
   U5657 : MUX2_X1 port map( A => REGISTERS_25_57_port, B => n5817, S => n37, Z
                           => n2897);
   U5658 : MUX2_X1 port map( A => REGISTERS_25_56_port, B => n5818, S => n37, Z
                           => n2896);
   U5659 : MUX2_X1 port map( A => REGISTERS_25_55_port, B => n5819, S => n37, Z
                           => n2895);
   U5660 : MUX2_X1 port map( A => REGISTERS_25_54_port, B => n5820, S => n37, Z
                           => n2894);
   U5661 : MUX2_X1 port map( A => REGISTERS_25_53_port, B => n5821, S => n37, Z
                           => n2893);
   U5662 : MUX2_X1 port map( A => REGISTERS_25_52_port, B => n5822, S => n37, Z
                           => n2892);
   U5663 : MUX2_X1 port map( A => REGISTERS_25_51_port, B => n5823, S => n37, Z
                           => n2891);
   U5664 : MUX2_X1 port map( A => REGISTERS_25_50_port, B => n5824, S => n37, Z
                           => n2890);
   U5665 : MUX2_X1 port map( A => REGISTERS_25_49_port, B => n5825, S => n37, Z
                           => n2889);
   U5666 : MUX2_X1 port map( A => REGISTERS_25_48_port, B => n5826, S => n37, Z
                           => n2888);
   U5667 : MUX2_X1 port map( A => REGISTERS_25_47_port, B => n5827, S => n37, Z
                           => n2887);
   U5668 : MUX2_X1 port map( A => REGISTERS_25_46_port, B => n5828, S => n37, Z
                           => n2886);
   U5669 : MUX2_X1 port map( A => REGISTERS_25_45_port, B => n5829, S => n37, Z
                           => n2885);
   U5670 : MUX2_X1 port map( A => REGISTERS_25_44_port, B => n5830, S => n37, Z
                           => n2884);
   U5671 : MUX2_X1 port map( A => REGISTERS_25_43_port, B => n5831, S => n37, Z
                           => n2883);
   U5672 : MUX2_X1 port map( A => REGISTERS_25_42_port, B => n5832, S => n37, Z
                           => n2882);
   U5673 : MUX2_X1 port map( A => REGISTERS_25_41_port, B => n5833, S => n37, Z
                           => n2881);
   U5674 : MUX2_X1 port map( A => REGISTERS_25_40_port, B => n5834, S => n37, Z
                           => n2880);
   U5675 : MUX2_X1 port map( A => REGISTERS_25_39_port, B => n5835, S => n37, Z
                           => n2879);
   U5676 : MUX2_X1 port map( A => REGISTERS_25_38_port, B => n5836, S => n37, Z
                           => n2878);
   U5677 : MUX2_X1 port map( A => REGISTERS_25_37_port, B => n5837, S => n37, Z
                           => n2877);
   U5678 : MUX2_X1 port map( A => REGISTERS_25_36_port, B => n5838, S => n37, Z
                           => n2876);
   U5679 : MUX2_X1 port map( A => REGISTERS_25_35_port, B => n5839, S => n37, Z
                           => n2875);
   U5680 : MUX2_X1 port map( A => REGISTERS_25_34_port, B => n5840, S => n37, Z
                           => n2874);
   U5681 : MUX2_X1 port map( A => REGISTERS_25_33_port, B => n5841, S => n37, Z
                           => n2873);
   U5682 : MUX2_X1 port map( A => REGISTERS_25_32_port, B => n5842, S => n37, Z
                           => n2872);
   U5683 : MUX2_X1 port map( A => REGISTERS_25_31_port, B => n5843, S => n37, Z
                           => n2871);
   U5684 : MUX2_X1 port map( A => REGISTERS_25_30_port, B => n5844, S => n37, Z
                           => n2870);
   U5685 : MUX2_X1 port map( A => REGISTERS_25_29_port, B => n5845, S => n37, Z
                           => n2869);
   U5686 : MUX2_X1 port map( A => REGISTERS_25_28_port, B => n5846, S => n37, Z
                           => n2868);
   U5687 : MUX2_X1 port map( A => REGISTERS_25_27_port, B => n5847, S => n37, Z
                           => n2867);
   U5688 : MUX2_X1 port map( A => REGISTERS_25_26_port, B => n5848, S => n37, Z
                           => n2866);
   U5689 : MUX2_X1 port map( A => REGISTERS_25_25_port, B => n5849, S => n37, Z
                           => n2865);
   U5690 : MUX2_X1 port map( A => REGISTERS_25_24_port, B => n5850, S => n37, Z
                           => n2864);
   U5691 : MUX2_X1 port map( A => REGISTERS_25_23_port, B => n5851, S => n37, Z
                           => n2863);
   U5692 : MUX2_X1 port map( A => REGISTERS_25_22_port, B => n5852, S => n37, Z
                           => n2862);
   U5693 : MUX2_X1 port map( A => REGISTERS_25_21_port, B => n5853, S => n37, Z
                           => n2861);
   U5694 : MUX2_X1 port map( A => REGISTERS_25_20_port, B => n5854, S => n37, Z
                           => n2860);
   U5695 : MUX2_X1 port map( A => REGISTERS_25_19_port, B => n5855, S => n37, Z
                           => n2859);
   U5696 : MUX2_X1 port map( A => REGISTERS_25_18_port, B => n5856, S => n37, Z
                           => n2858);
   U5697 : MUX2_X1 port map( A => REGISTERS_25_17_port, B => n5857, S => n37, Z
                           => n2857);
   U5698 : MUX2_X1 port map( A => REGISTERS_25_16_port, B => n5858, S => n37, Z
                           => n2856);
   U5699 : MUX2_X1 port map( A => REGISTERS_25_15_port, B => n5859, S => n37, Z
                           => n2855);
   U5700 : MUX2_X1 port map( A => REGISTERS_25_14_port, B => n5860, S => n37, Z
                           => n2854);
   U5701 : MUX2_X1 port map( A => REGISTERS_25_13_port, B => n5861, S => n37, Z
                           => n2853);
   U5702 : MUX2_X1 port map( A => REGISTERS_25_12_port, B => n5862, S => n37, Z
                           => n2852);
   U5703 : MUX2_X1 port map( A => REGISTERS_25_11_port, B => n5863, S => n37, Z
                           => n2851);
   U5704 : MUX2_X1 port map( A => REGISTERS_25_10_port, B => n5864, S => n37, Z
                           => n2850);
   U5705 : MUX2_X1 port map( A => REGISTERS_25_9_port, B => n5865, S => n37, Z 
                           => n2849);
   U5706 : MUX2_X1 port map( A => REGISTERS_25_8_port, B => n5866, S => n37, Z 
                           => n2848);
   U5707 : MUX2_X1 port map( A => REGISTERS_25_7_port, B => n5867, S => n37, Z 
                           => n2847);
   U5708 : MUX2_X1 port map( A => REGISTERS_25_6_port, B => n5868, S => n37, Z 
                           => n2846);
   U5709 : MUX2_X1 port map( A => REGISTERS_25_5_port, B => n5869, S => n37, Z 
                           => n2845);
   U5710 : MUX2_X1 port map( A => REGISTERS_25_4_port, B => n5870, S => n37, Z 
                           => n2844);
   U5711 : MUX2_X1 port map( A => REGISTERS_25_3_port, B => n5871, S => n37, Z 
                           => n2843);
   U5712 : MUX2_X1 port map( A => REGISTERS_25_2_port, B => n5872, S => n37, Z 
                           => n2842);
   U5713 : MUX2_X1 port map( A => REGISTERS_25_1_port, B => n5873, S => n37, Z 
                           => n2841);
   U5714 : MUX2_X1 port map( A => REGISTERS_25_0_port, B => n5874, S => n37, Z 
                           => n2840);
   U5715 : OAI21_X1 port map( B1 => n5878, B2 => n5913, A => n5744, ZN => n5917
                           );
   U5716 : NAND3_X1 port map( A1 => n5914, A2 => n5915, A3 => ADD_WR(0), ZN => 
                           n5878);
   U5717 : MUX2_X1 port map( A => REGISTERS_26_63_port, B => n5810, S => n39, Z
                           => n2839);
   U5718 : MUX2_X1 port map( A => REGISTERS_26_62_port, B => n5812, S => n39, Z
                           => n2838);
   U5719 : MUX2_X1 port map( A => REGISTERS_26_61_port, B => n5813, S => n39, Z
                           => n2837);
   U5720 : MUX2_X1 port map( A => REGISTERS_26_60_port, B => n5814, S => n39, Z
                           => n2836);
   U5721 : MUX2_X1 port map( A => REGISTERS_26_59_port, B => n5815, S => n39, Z
                           => n2835);
   U5722 : MUX2_X1 port map( A => REGISTERS_26_58_port, B => n5816, S => n39, Z
                           => n2834);
   U5723 : MUX2_X1 port map( A => REGISTERS_26_57_port, B => n5817, S => n39, Z
                           => n2833);
   U5724 : MUX2_X1 port map( A => REGISTERS_26_56_port, B => n5818, S => n39, Z
                           => n2832);
   U5725 : MUX2_X1 port map( A => REGISTERS_26_55_port, B => n5819, S => n39, Z
                           => n2831);
   U5726 : MUX2_X1 port map( A => REGISTERS_26_54_port, B => n5820, S => n39, Z
                           => n2830);
   U5727 : MUX2_X1 port map( A => REGISTERS_26_53_port, B => n5821, S => n39, Z
                           => n2829);
   U5728 : MUX2_X1 port map( A => REGISTERS_26_52_port, B => n5822, S => n39, Z
                           => n2828);
   U5729 : MUX2_X1 port map( A => REGISTERS_26_51_port, B => n5823, S => n39, Z
                           => n2827);
   U5730 : MUX2_X1 port map( A => REGISTERS_26_50_port, B => n5824, S => n39, Z
                           => n2826);
   U5731 : MUX2_X1 port map( A => REGISTERS_26_49_port, B => n5825, S => n39, Z
                           => n2825);
   U5732 : MUX2_X1 port map( A => REGISTERS_26_48_port, B => n5826, S => n39, Z
                           => n2824);
   U5733 : MUX2_X1 port map( A => REGISTERS_26_47_port, B => n5827, S => n39, Z
                           => n2823);
   U5734 : MUX2_X1 port map( A => REGISTERS_26_46_port, B => n5828, S => n39, Z
                           => n2822);
   U5735 : MUX2_X1 port map( A => REGISTERS_26_45_port, B => n5829, S => n39, Z
                           => n2821);
   U5736 : MUX2_X1 port map( A => REGISTERS_26_44_port, B => n5830, S => n39, Z
                           => n2820);
   U5737 : MUX2_X1 port map( A => REGISTERS_26_43_port, B => n5831, S => n39, Z
                           => n2819);
   U5738 : MUX2_X1 port map( A => REGISTERS_26_42_port, B => n5832, S => n39, Z
                           => n2818);
   U5739 : MUX2_X1 port map( A => REGISTERS_26_41_port, B => n5833, S => n39, Z
                           => n2817);
   U5740 : MUX2_X1 port map( A => REGISTERS_26_40_port, B => n5834, S => n39, Z
                           => n2816);
   U5741 : MUX2_X1 port map( A => REGISTERS_26_39_port, B => n5835, S => n39, Z
                           => n2815);
   U5742 : MUX2_X1 port map( A => REGISTERS_26_38_port, B => n5836, S => n39, Z
                           => n2814);
   U5743 : MUX2_X1 port map( A => REGISTERS_26_37_port, B => n5837, S => n39, Z
                           => n2813);
   U5744 : MUX2_X1 port map( A => REGISTERS_26_36_port, B => n5838, S => n39, Z
                           => n2812);
   U5745 : MUX2_X1 port map( A => REGISTERS_26_35_port, B => n5839, S => n39, Z
                           => n2811);
   U5746 : MUX2_X1 port map( A => REGISTERS_26_34_port, B => n5840, S => n39, Z
                           => n2810);
   U5747 : MUX2_X1 port map( A => REGISTERS_26_33_port, B => n5841, S => n39, Z
                           => n2809);
   U5748 : MUX2_X1 port map( A => REGISTERS_26_32_port, B => n5842, S => n39, Z
                           => n2808);
   U5749 : MUX2_X1 port map( A => REGISTERS_26_31_port, B => n5843, S => n39, Z
                           => n2807);
   U5750 : MUX2_X1 port map( A => REGISTERS_26_30_port, B => n5844, S => n39, Z
                           => n2806);
   U5751 : MUX2_X1 port map( A => REGISTERS_26_29_port, B => n5845, S => n39, Z
                           => n2805);
   U5752 : MUX2_X1 port map( A => REGISTERS_26_28_port, B => n5846, S => n39, Z
                           => n2804);
   U5753 : MUX2_X1 port map( A => REGISTERS_26_27_port, B => n5847, S => n39, Z
                           => n2803);
   U5754 : MUX2_X1 port map( A => REGISTERS_26_26_port, B => n5848, S => n39, Z
                           => n2802);
   U5755 : MUX2_X1 port map( A => REGISTERS_26_25_port, B => n5849, S => n39, Z
                           => n2801);
   U5756 : MUX2_X1 port map( A => REGISTERS_26_24_port, B => n5850, S => n39, Z
                           => n2800);
   U5757 : MUX2_X1 port map( A => REGISTERS_26_23_port, B => n5851, S => n39, Z
                           => n2799);
   U5758 : MUX2_X1 port map( A => REGISTERS_26_22_port, B => n5852, S => n39, Z
                           => n2798);
   U5759 : MUX2_X1 port map( A => REGISTERS_26_21_port, B => n5853, S => n39, Z
                           => n2797);
   U5760 : MUX2_X1 port map( A => REGISTERS_26_20_port, B => n5854, S => n39, Z
                           => n2796);
   U5761 : MUX2_X1 port map( A => REGISTERS_26_19_port, B => n5855, S => n39, Z
                           => n2795);
   U5762 : MUX2_X1 port map( A => REGISTERS_26_18_port, B => n5856, S => n39, Z
                           => n2794);
   U5763 : MUX2_X1 port map( A => REGISTERS_26_17_port, B => n5857, S => n39, Z
                           => n2793);
   U5764 : MUX2_X1 port map( A => REGISTERS_26_16_port, B => n5858, S => n39, Z
                           => n2792);
   U5765 : MUX2_X1 port map( A => REGISTERS_26_15_port, B => n5859, S => n39, Z
                           => n2791);
   U5766 : MUX2_X1 port map( A => REGISTERS_26_14_port, B => n5860, S => n39, Z
                           => n2790);
   U5767 : MUX2_X1 port map( A => REGISTERS_26_13_port, B => n5861, S => n39, Z
                           => n2789);
   U5768 : MUX2_X1 port map( A => REGISTERS_26_12_port, B => n5862, S => n39, Z
                           => n2788);
   U5769 : MUX2_X1 port map( A => REGISTERS_26_11_port, B => n5863, S => n39, Z
                           => n2787);
   U5770 : MUX2_X1 port map( A => REGISTERS_26_10_port, B => n5864, S => n39, Z
                           => n2786);
   U5771 : MUX2_X1 port map( A => REGISTERS_26_9_port, B => n5865, S => n39, Z 
                           => n2785);
   U5772 : MUX2_X1 port map( A => REGISTERS_26_8_port, B => n5866, S => n39, Z 
                           => n2784);
   U5773 : MUX2_X1 port map( A => REGISTERS_26_7_port, B => n5867, S => n39, Z 
                           => n2783);
   U5774 : MUX2_X1 port map( A => REGISTERS_26_6_port, B => n5868, S => n39, Z 
                           => n2782);
   U5775 : MUX2_X1 port map( A => REGISTERS_26_5_port, B => n5869, S => n39, Z 
                           => n2781);
   U5776 : MUX2_X1 port map( A => REGISTERS_26_4_port, B => n5870, S => n39, Z 
                           => n2780);
   U5777 : MUX2_X1 port map( A => REGISTERS_26_3_port, B => n5871, S => n39, Z 
                           => n2779);
   U5778 : MUX2_X1 port map( A => REGISTERS_26_2_port, B => n5872, S => n39, Z 
                           => n2778);
   U5779 : MUX2_X1 port map( A => REGISTERS_26_1_port, B => n5873, S => n39, Z 
                           => n2777);
   U5780 : MUX2_X1 port map( A => REGISTERS_26_0_port, B => n5874, S => n39, Z 
                           => n2776);
   U5781 : OAI21_X1 port map( B1 => n5880, B2 => n5913, A => n5744, ZN => n5918
                           );
   U5782 : NAND3_X1 port map( A1 => n5916, A2 => n5915, A3 => ADD_WR(1), ZN => 
                           n5880);
   U5783 : MUX2_X1 port map( A => REGISTERS_27_63_port, B => n5810, S => n33, Z
                           => n2775);
   U5784 : MUX2_X1 port map( A => REGISTERS_27_62_port, B => n5812, S => n33, Z
                           => n2774);
   U5785 : MUX2_X1 port map( A => REGISTERS_27_61_port, B => n5813, S => n33, Z
                           => n2773);
   U5786 : MUX2_X1 port map( A => REGISTERS_27_60_port, B => n5814, S => n33, Z
                           => n2772);
   U5787 : MUX2_X1 port map( A => REGISTERS_27_59_port, B => n5815, S => n33, Z
                           => n2771);
   U5788 : MUX2_X1 port map( A => REGISTERS_27_58_port, B => n5816, S => n33, Z
                           => n2770);
   U5789 : MUX2_X1 port map( A => REGISTERS_27_57_port, B => n5817, S => n33, Z
                           => n2769);
   U5790 : MUX2_X1 port map( A => REGISTERS_27_56_port, B => n5818, S => n33, Z
                           => n2768);
   U5791 : MUX2_X1 port map( A => REGISTERS_27_55_port, B => n5819, S => n33, Z
                           => n2767);
   U5792 : MUX2_X1 port map( A => REGISTERS_27_54_port, B => n5820, S => n33, Z
                           => n2766);
   U5793 : MUX2_X1 port map( A => REGISTERS_27_53_port, B => n5821, S => n33, Z
                           => n2765);
   U5794 : MUX2_X1 port map( A => REGISTERS_27_52_port, B => n5822, S => n33, Z
                           => n2764);
   U5795 : MUX2_X1 port map( A => REGISTERS_27_51_port, B => n5823, S => n33, Z
                           => n2763);
   U5796 : MUX2_X1 port map( A => REGISTERS_27_50_port, B => n5824, S => n33, Z
                           => n2762);
   U5797 : MUX2_X1 port map( A => REGISTERS_27_49_port, B => n5825, S => n33, Z
                           => n2761);
   U5798 : MUX2_X1 port map( A => REGISTERS_27_48_port, B => n5826, S => n33, Z
                           => n2760);
   U5799 : MUX2_X1 port map( A => REGISTERS_27_47_port, B => n5827, S => n33, Z
                           => n2759);
   U5800 : MUX2_X1 port map( A => REGISTERS_27_46_port, B => n5828, S => n33, Z
                           => n2758);
   U5801 : MUX2_X1 port map( A => REGISTERS_27_45_port, B => n5829, S => n33, Z
                           => n2757);
   U5802 : MUX2_X1 port map( A => REGISTERS_27_44_port, B => n5830, S => n33, Z
                           => n2756);
   U5803 : MUX2_X1 port map( A => REGISTERS_27_43_port, B => n5831, S => n33, Z
                           => n2755);
   U5804 : MUX2_X1 port map( A => REGISTERS_27_42_port, B => n5832, S => n33, Z
                           => n2754);
   U5805 : MUX2_X1 port map( A => REGISTERS_27_41_port, B => n5833, S => n33, Z
                           => n2753);
   U5806 : MUX2_X1 port map( A => REGISTERS_27_40_port, B => n5834, S => n33, Z
                           => n2752);
   U5807 : MUX2_X1 port map( A => REGISTERS_27_39_port, B => n5835, S => n33, Z
                           => n2751);
   U5808 : MUX2_X1 port map( A => REGISTERS_27_38_port, B => n5836, S => n33, Z
                           => n2750);
   U5809 : MUX2_X1 port map( A => REGISTERS_27_37_port, B => n5837, S => n33, Z
                           => n2749);
   U5810 : MUX2_X1 port map( A => REGISTERS_27_36_port, B => n5838, S => n33, Z
                           => n2748);
   U5811 : MUX2_X1 port map( A => REGISTERS_27_35_port, B => n5839, S => n33, Z
                           => n2747);
   U5812 : MUX2_X1 port map( A => REGISTERS_27_34_port, B => n5840, S => n33, Z
                           => n2746);
   U5813 : MUX2_X1 port map( A => REGISTERS_27_33_port, B => n5841, S => n33, Z
                           => n2745);
   U5814 : MUX2_X1 port map( A => REGISTERS_27_32_port, B => n5842, S => n33, Z
                           => n2744);
   U5815 : MUX2_X1 port map( A => REGISTERS_27_31_port, B => n5843, S => n33, Z
                           => n2743);
   U5816 : MUX2_X1 port map( A => REGISTERS_27_30_port, B => n5844, S => n33, Z
                           => n2742);
   U5817 : MUX2_X1 port map( A => REGISTERS_27_29_port, B => n5845, S => n33, Z
                           => n2741);
   U5818 : MUX2_X1 port map( A => REGISTERS_27_28_port, B => n5846, S => n33, Z
                           => n2740);
   U5819 : MUX2_X1 port map( A => REGISTERS_27_27_port, B => n5847, S => n33, Z
                           => n2739);
   U5820 : MUX2_X1 port map( A => REGISTERS_27_26_port, B => n5848, S => n33, Z
                           => n2738);
   U5821 : MUX2_X1 port map( A => REGISTERS_27_25_port, B => n5849, S => n33, Z
                           => n2737);
   U5822 : MUX2_X1 port map( A => REGISTERS_27_24_port, B => n5850, S => n33, Z
                           => n2736);
   U5823 : MUX2_X1 port map( A => REGISTERS_27_23_port, B => n5851, S => n33, Z
                           => n2735);
   U5824 : MUX2_X1 port map( A => REGISTERS_27_22_port, B => n5852, S => n33, Z
                           => n2734);
   U5825 : MUX2_X1 port map( A => REGISTERS_27_21_port, B => n5853, S => n33, Z
                           => n2733);
   U5826 : MUX2_X1 port map( A => REGISTERS_27_20_port, B => n5854, S => n33, Z
                           => n2732);
   U5827 : MUX2_X1 port map( A => REGISTERS_27_19_port, B => n5855, S => n33, Z
                           => n2731);
   U5828 : MUX2_X1 port map( A => REGISTERS_27_18_port, B => n5856, S => n33, Z
                           => n2730);
   U5829 : MUX2_X1 port map( A => REGISTERS_27_17_port, B => n5857, S => n33, Z
                           => n2729);
   U5830 : MUX2_X1 port map( A => REGISTERS_27_16_port, B => n5858, S => n33, Z
                           => n2728);
   U5831 : MUX2_X1 port map( A => REGISTERS_27_15_port, B => n5859, S => n33, Z
                           => n2727);
   U5832 : MUX2_X1 port map( A => REGISTERS_27_14_port, B => n5860, S => n33, Z
                           => n2726);
   U5833 : MUX2_X1 port map( A => REGISTERS_27_13_port, B => n5861, S => n33, Z
                           => n2725);
   U5834 : MUX2_X1 port map( A => REGISTERS_27_12_port, B => n5862, S => n33, Z
                           => n2724);
   U5835 : MUX2_X1 port map( A => REGISTERS_27_11_port, B => n5863, S => n33, Z
                           => n2723);
   U5836 : MUX2_X1 port map( A => REGISTERS_27_10_port, B => n5864, S => n33, Z
                           => n2722);
   U5837 : MUX2_X1 port map( A => REGISTERS_27_9_port, B => n5865, S => n33, Z 
                           => n2721);
   U5838 : MUX2_X1 port map( A => REGISTERS_27_8_port, B => n5866, S => n33, Z 
                           => n2720);
   U5839 : MUX2_X1 port map( A => REGISTERS_27_7_port, B => n5867, S => n33, Z 
                           => n2719);
   U5840 : MUX2_X1 port map( A => REGISTERS_27_6_port, B => n5868, S => n33, Z 
                           => n2718);
   U5841 : MUX2_X1 port map( A => REGISTERS_27_5_port, B => n5869, S => n33, Z 
                           => n2717);
   U5842 : MUX2_X1 port map( A => REGISTERS_27_4_port, B => n5870, S => n33, Z 
                           => n2716);
   U5843 : MUX2_X1 port map( A => REGISTERS_27_3_port, B => n5871, S => n33, Z 
                           => n2715);
   U5844 : MUX2_X1 port map( A => REGISTERS_27_2_port, B => n5872, S => n33, Z 
                           => n2714);
   U5845 : MUX2_X1 port map( A => REGISTERS_27_1_port, B => n5873, S => n33, Z 
                           => n2713);
   U5846 : MUX2_X1 port map( A => REGISTERS_27_0_port, B => n5874, S => n33, Z 
                           => n2712);
   U5847 : OAI21_X1 port map( B1 => n5882, B2 => n5913, A => n5744, ZN => n5919
                           );
   U5848 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n5915, A3 => ADD_WR(1), ZN
                           => n5882);
   U5849 : INV_X1 port map( A => ADD_WR(2), ZN => n5915);
   U5850 : MUX2_X1 port map( A => REGISTERS_28_63_port, B => n5810, S => n35, Z
                           => n2711);
   U5851 : MUX2_X1 port map( A => REGISTERS_28_62_port, B => n5812, S => n35, Z
                           => n2710);
   U5852 : MUX2_X1 port map( A => REGISTERS_28_61_port, B => n5813, S => n35, Z
                           => n2709);
   U5853 : MUX2_X1 port map( A => REGISTERS_28_60_port, B => n5814, S => n35, Z
                           => n2708);
   U5854 : MUX2_X1 port map( A => REGISTERS_28_59_port, B => n5815, S => n35, Z
                           => n2707);
   U5855 : MUX2_X1 port map( A => REGISTERS_28_58_port, B => n5816, S => n35, Z
                           => n2706);
   U5856 : MUX2_X1 port map( A => REGISTERS_28_57_port, B => n5817, S => n35, Z
                           => n2705);
   U5857 : MUX2_X1 port map( A => REGISTERS_28_56_port, B => n5818, S => n35, Z
                           => n2704);
   U5858 : MUX2_X1 port map( A => REGISTERS_28_55_port, B => n5819, S => n35, Z
                           => n2703);
   U5859 : MUX2_X1 port map( A => REGISTERS_28_54_port, B => n5820, S => n35, Z
                           => n2702);
   U5860 : MUX2_X1 port map( A => REGISTERS_28_53_port, B => n5821, S => n35, Z
                           => n2701);
   U5861 : MUX2_X1 port map( A => REGISTERS_28_52_port, B => n5822, S => n35, Z
                           => n2700);
   U5862 : MUX2_X1 port map( A => REGISTERS_28_51_port, B => n5823, S => n35, Z
                           => n2699);
   U5863 : MUX2_X1 port map( A => REGISTERS_28_50_port, B => n5824, S => n35, Z
                           => n2698);
   U5864 : MUX2_X1 port map( A => REGISTERS_28_49_port, B => n5825, S => n35, Z
                           => n2697);
   U5865 : MUX2_X1 port map( A => REGISTERS_28_48_port, B => n5826, S => n35, Z
                           => n2696);
   U5866 : MUX2_X1 port map( A => REGISTERS_28_47_port, B => n5827, S => n35, Z
                           => n2695);
   U5867 : MUX2_X1 port map( A => REGISTERS_28_46_port, B => n5828, S => n35, Z
                           => n2694);
   U5868 : MUX2_X1 port map( A => REGISTERS_28_45_port, B => n5829, S => n35, Z
                           => n2693);
   U5869 : MUX2_X1 port map( A => REGISTERS_28_44_port, B => n5830, S => n35, Z
                           => n2692);
   U5870 : MUX2_X1 port map( A => REGISTERS_28_43_port, B => n5831, S => n35, Z
                           => n2691);
   U5871 : MUX2_X1 port map( A => REGISTERS_28_42_port, B => n5832, S => n35, Z
                           => n2690);
   U5872 : MUX2_X1 port map( A => REGISTERS_28_41_port, B => n5833, S => n35, Z
                           => n2689);
   U5873 : MUX2_X1 port map( A => REGISTERS_28_40_port, B => n5834, S => n35, Z
                           => n2688);
   U5874 : MUX2_X1 port map( A => REGISTERS_28_39_port, B => n5835, S => n35, Z
                           => n2687);
   U5875 : MUX2_X1 port map( A => REGISTERS_28_38_port, B => n5836, S => n35, Z
                           => n2686);
   U5876 : MUX2_X1 port map( A => REGISTERS_28_37_port, B => n5837, S => n35, Z
                           => n2685);
   U5877 : MUX2_X1 port map( A => REGISTERS_28_36_port, B => n5838, S => n35, Z
                           => n2684);
   U5878 : MUX2_X1 port map( A => REGISTERS_28_35_port, B => n5839, S => n35, Z
                           => n2683);
   U5879 : MUX2_X1 port map( A => REGISTERS_28_34_port, B => n5840, S => n35, Z
                           => n2682);
   U5880 : MUX2_X1 port map( A => REGISTERS_28_33_port, B => n5841, S => n35, Z
                           => n2681);
   U5881 : MUX2_X1 port map( A => REGISTERS_28_32_port, B => n5842, S => n35, Z
                           => n2680);
   U5882 : MUX2_X1 port map( A => REGISTERS_28_31_port, B => n5843, S => n35, Z
                           => n2679);
   U5883 : MUX2_X1 port map( A => REGISTERS_28_30_port, B => n5844, S => n35, Z
                           => n2678);
   U5884 : MUX2_X1 port map( A => REGISTERS_28_29_port, B => n5845, S => n35, Z
                           => n2677);
   U5885 : MUX2_X1 port map( A => REGISTERS_28_28_port, B => n5846, S => n35, Z
                           => n2676);
   U5886 : MUX2_X1 port map( A => REGISTERS_28_27_port, B => n5847, S => n35, Z
                           => n2675);
   U5887 : MUX2_X1 port map( A => REGISTERS_28_26_port, B => n5848, S => n35, Z
                           => n2674);
   U5888 : MUX2_X1 port map( A => REGISTERS_28_25_port, B => n5849, S => n35, Z
                           => n2673);
   U5889 : MUX2_X1 port map( A => REGISTERS_28_24_port, B => n5850, S => n35, Z
                           => n2672);
   U5890 : MUX2_X1 port map( A => REGISTERS_28_23_port, B => n5851, S => n35, Z
                           => n2671);
   U5891 : MUX2_X1 port map( A => REGISTERS_28_22_port, B => n5852, S => n35, Z
                           => n2670);
   U5892 : MUX2_X1 port map( A => REGISTERS_28_21_port, B => n5853, S => n35, Z
                           => n2669);
   U5893 : MUX2_X1 port map( A => REGISTERS_28_20_port, B => n5854, S => n35, Z
                           => n2668);
   U5894 : MUX2_X1 port map( A => REGISTERS_28_19_port, B => n5855, S => n35, Z
                           => n2667);
   U5895 : MUX2_X1 port map( A => REGISTERS_28_18_port, B => n5856, S => n35, Z
                           => n2666);
   U5896 : MUX2_X1 port map( A => REGISTERS_28_17_port, B => n5857, S => n35, Z
                           => n2665);
   U5897 : MUX2_X1 port map( A => REGISTERS_28_16_port, B => n5858, S => n35, Z
                           => n2664);
   U5898 : MUX2_X1 port map( A => REGISTERS_28_15_port, B => n5859, S => n35, Z
                           => n2663);
   U5899 : MUX2_X1 port map( A => REGISTERS_28_14_port, B => n5860, S => n35, Z
                           => n2662);
   U5900 : MUX2_X1 port map( A => REGISTERS_28_13_port, B => n5861, S => n35, Z
                           => n2661);
   U5901 : MUX2_X1 port map( A => REGISTERS_28_12_port, B => n5862, S => n35, Z
                           => n2660);
   U5902 : MUX2_X1 port map( A => REGISTERS_28_11_port, B => n5863, S => n35, Z
                           => n2659);
   U5903 : MUX2_X1 port map( A => REGISTERS_28_10_port, B => n5864, S => n35, Z
                           => n2658);
   U5904 : MUX2_X1 port map( A => REGISTERS_28_9_port, B => n5865, S => n35, Z 
                           => n2657);
   U5905 : MUX2_X1 port map( A => REGISTERS_28_8_port, B => n5866, S => n35, Z 
                           => n2656);
   U5906 : MUX2_X1 port map( A => REGISTERS_28_7_port, B => n5867, S => n35, Z 
                           => n2655);
   U5907 : MUX2_X1 port map( A => REGISTERS_28_6_port, B => n5868, S => n35, Z 
                           => n2654);
   U5908 : MUX2_X1 port map( A => REGISTERS_28_5_port, B => n5869, S => n35, Z 
                           => n2653);
   U5909 : MUX2_X1 port map( A => REGISTERS_28_4_port, B => n5870, S => n35, Z 
                           => n2652);
   U5910 : MUX2_X1 port map( A => REGISTERS_28_3_port, B => n5871, S => n35, Z 
                           => n2651);
   U5911 : MUX2_X1 port map( A => REGISTERS_28_2_port, B => n5872, S => n35, Z 
                           => n2650);
   U5912 : MUX2_X1 port map( A => REGISTERS_28_1_port, B => n5873, S => n35, Z 
                           => n2649);
   U5913 : MUX2_X1 port map( A => REGISTERS_28_0_port, B => n5874, S => n35, Z 
                           => n2648);
   U5914 : OAI21_X1 port map( B1 => n5884, B2 => n5913, A => n5744, ZN => n5920
                           );
   U5915 : NAND3_X1 port map( A1 => n5916, A2 => n5914, A3 => ADD_WR(2), ZN => 
                           n5884);
   U5916 : MUX2_X1 port map( A => REGISTERS_29_63_port, B => n5810, S => n29, Z
                           => n2647);
   U5917 : MUX2_X1 port map( A => REGISTERS_29_62_port, B => n5812, S => n29, Z
                           => n2646);
   U5918 : MUX2_X1 port map( A => REGISTERS_29_61_port, B => n5813, S => n29, Z
                           => n2645);
   U5919 : MUX2_X1 port map( A => REGISTERS_29_60_port, B => n5814, S => n29, Z
                           => n2644);
   U5920 : MUX2_X1 port map( A => REGISTERS_29_59_port, B => n5815, S => n29, Z
                           => n2643);
   U5921 : MUX2_X1 port map( A => REGISTERS_29_58_port, B => n5816, S => n29, Z
                           => n2642);
   U5922 : MUX2_X1 port map( A => REGISTERS_29_57_port, B => n5817, S => n29, Z
                           => n2641);
   U5923 : MUX2_X1 port map( A => REGISTERS_29_56_port, B => n5818, S => n29, Z
                           => n2640);
   U5924 : MUX2_X1 port map( A => REGISTERS_29_55_port, B => n5819, S => n29, Z
                           => n2639);
   U5925 : MUX2_X1 port map( A => REGISTERS_29_54_port, B => n5820, S => n29, Z
                           => n2638);
   U5926 : MUX2_X1 port map( A => REGISTERS_29_53_port, B => n5821, S => n29, Z
                           => n2637);
   U5927 : MUX2_X1 port map( A => REGISTERS_29_52_port, B => n5822, S => n29, Z
                           => n2636);
   U5928 : MUX2_X1 port map( A => REGISTERS_29_51_port, B => n5823, S => n29, Z
                           => n2635);
   U5929 : MUX2_X1 port map( A => REGISTERS_29_50_port, B => n5824, S => n29, Z
                           => n2634);
   U5930 : MUX2_X1 port map( A => REGISTERS_29_49_port, B => n5825, S => n29, Z
                           => n2633);
   U5931 : MUX2_X1 port map( A => REGISTERS_29_48_port, B => n5826, S => n29, Z
                           => n2632);
   U5932 : MUX2_X1 port map( A => REGISTERS_29_47_port, B => n5827, S => n29, Z
                           => n2631);
   U5933 : MUX2_X1 port map( A => REGISTERS_29_46_port, B => n5828, S => n29, Z
                           => n2630);
   U5934 : MUX2_X1 port map( A => REGISTERS_29_45_port, B => n5829, S => n29, Z
                           => n2629);
   U5935 : MUX2_X1 port map( A => REGISTERS_29_44_port, B => n5830, S => n29, Z
                           => n2628);
   U5936 : MUX2_X1 port map( A => REGISTERS_29_43_port, B => n5831, S => n29, Z
                           => n2627);
   U5937 : MUX2_X1 port map( A => REGISTERS_29_42_port, B => n5832, S => n29, Z
                           => n2626);
   U5938 : MUX2_X1 port map( A => REGISTERS_29_41_port, B => n5833, S => n29, Z
                           => n2625);
   U5939 : MUX2_X1 port map( A => REGISTERS_29_40_port, B => n5834, S => n29, Z
                           => n2624);
   U5940 : MUX2_X1 port map( A => REGISTERS_29_39_port, B => n5835, S => n29, Z
                           => n2623);
   U5941 : MUX2_X1 port map( A => REGISTERS_29_38_port, B => n5836, S => n29, Z
                           => n2622);
   U5942 : MUX2_X1 port map( A => REGISTERS_29_37_port, B => n5837, S => n29, Z
                           => n2621);
   U5943 : MUX2_X1 port map( A => REGISTERS_29_36_port, B => n5838, S => n29, Z
                           => n2620);
   U5944 : MUX2_X1 port map( A => REGISTERS_29_35_port, B => n5839, S => n29, Z
                           => n2619);
   U5945 : MUX2_X1 port map( A => REGISTERS_29_34_port, B => n5840, S => n29, Z
                           => n2618);
   U5946 : MUX2_X1 port map( A => REGISTERS_29_33_port, B => n5841, S => n29, Z
                           => n2617);
   U5947 : MUX2_X1 port map( A => REGISTERS_29_32_port, B => n5842, S => n29, Z
                           => n2616);
   U5948 : MUX2_X1 port map( A => REGISTERS_29_31_port, B => n5843, S => n29, Z
                           => n2615);
   U5949 : MUX2_X1 port map( A => REGISTERS_29_30_port, B => n5844, S => n29, Z
                           => n2614);
   U5950 : MUX2_X1 port map( A => REGISTERS_29_29_port, B => n5845, S => n29, Z
                           => n2613);
   U5951 : MUX2_X1 port map( A => REGISTERS_29_28_port, B => n5846, S => n29, Z
                           => n2612);
   U5952 : MUX2_X1 port map( A => REGISTERS_29_27_port, B => n5847, S => n29, Z
                           => n2611);
   U5953 : MUX2_X1 port map( A => REGISTERS_29_26_port, B => n5848, S => n29, Z
                           => n2610);
   U5954 : MUX2_X1 port map( A => REGISTERS_29_25_port, B => n5849, S => n29, Z
                           => n2609);
   U5955 : MUX2_X1 port map( A => REGISTERS_29_24_port, B => n5850, S => n29, Z
                           => n2608);
   U5956 : MUX2_X1 port map( A => REGISTERS_29_23_port, B => n5851, S => n29, Z
                           => n2607);
   U5957 : MUX2_X1 port map( A => REGISTERS_29_22_port, B => n5852, S => n29, Z
                           => n2606);
   U5958 : MUX2_X1 port map( A => REGISTERS_29_21_port, B => n5853, S => n29, Z
                           => n2605);
   U5959 : MUX2_X1 port map( A => REGISTERS_29_20_port, B => n5854, S => n29, Z
                           => n2604);
   U5960 : MUX2_X1 port map( A => REGISTERS_29_19_port, B => n5855, S => n29, Z
                           => n2603);
   U5961 : MUX2_X1 port map( A => REGISTERS_29_18_port, B => n5856, S => n29, Z
                           => n2602);
   U5962 : MUX2_X1 port map( A => REGISTERS_29_17_port, B => n5857, S => n29, Z
                           => n2601);
   U5963 : MUX2_X1 port map( A => REGISTERS_29_16_port, B => n5858, S => n29, Z
                           => n2600);
   U5964 : MUX2_X1 port map( A => REGISTERS_29_15_port, B => n5859, S => n29, Z
                           => n2599);
   U5965 : MUX2_X1 port map( A => REGISTERS_29_14_port, B => n5860, S => n29, Z
                           => n2598);
   U5966 : MUX2_X1 port map( A => REGISTERS_29_13_port, B => n5861, S => n29, Z
                           => n2597);
   U5967 : MUX2_X1 port map( A => REGISTERS_29_12_port, B => n5862, S => n29, Z
                           => n2596);
   U5968 : MUX2_X1 port map( A => REGISTERS_29_11_port, B => n5863, S => n29, Z
                           => n2595);
   U5969 : MUX2_X1 port map( A => REGISTERS_29_10_port, B => n5864, S => n29, Z
                           => n2594);
   U5970 : MUX2_X1 port map( A => REGISTERS_29_9_port, B => n5865, S => n29, Z 
                           => n2593);
   U5971 : MUX2_X1 port map( A => REGISTERS_29_8_port, B => n5866, S => n29, Z 
                           => n2592);
   U5972 : MUX2_X1 port map( A => REGISTERS_29_7_port, B => n5867, S => n29, Z 
                           => n2591);
   U5973 : MUX2_X1 port map( A => REGISTERS_29_6_port, B => n5868, S => n29, Z 
                           => n2590);
   U5974 : MUX2_X1 port map( A => REGISTERS_29_5_port, B => n5869, S => n29, Z 
                           => n2589);
   U5975 : MUX2_X1 port map( A => REGISTERS_29_4_port, B => n5870, S => n29, Z 
                           => n2588);
   U5976 : MUX2_X1 port map( A => REGISTERS_29_3_port, B => n5871, S => n29, Z 
                           => n2587);
   U5977 : MUX2_X1 port map( A => REGISTERS_29_2_port, B => n5872, S => n29, Z 
                           => n2586);
   U5978 : MUX2_X1 port map( A => REGISTERS_29_1_port, B => n5873, S => n29, Z 
                           => n2585);
   U5979 : MUX2_X1 port map( A => REGISTERS_29_0_port, B => n5874, S => n29, Z 
                           => n2584);
   U5980 : OAI21_X1 port map( B1 => n5886, B2 => n5913, A => n5744, ZN => n5921
                           );
   U5981 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n5914, A3 => ADD_WR(2), ZN
                           => n5886);
   U5982 : INV_X1 port map( A => ADD_WR(1), ZN => n5914);
   U5983 : MUX2_X1 port map( A => REGISTERS_30_63_port, B => n5810, S => n31, Z
                           => n2583);
   U5984 : MUX2_X1 port map( A => REGISTERS_30_62_port, B => n5812, S => n31, Z
                           => n2582);
   U5985 : MUX2_X1 port map( A => REGISTERS_30_61_port, B => n5813, S => n31, Z
                           => n2581);
   U5986 : MUX2_X1 port map( A => REGISTERS_30_60_port, B => n5814, S => n31, Z
                           => n2580);
   U5987 : MUX2_X1 port map( A => REGISTERS_30_59_port, B => n5815, S => n31, Z
                           => n2579);
   U5988 : MUX2_X1 port map( A => REGISTERS_30_58_port, B => n5816, S => n31, Z
                           => n2578);
   U5989 : MUX2_X1 port map( A => REGISTERS_30_57_port, B => n5817, S => n31, Z
                           => n2577);
   U5990 : MUX2_X1 port map( A => REGISTERS_30_56_port, B => n5818, S => n31, Z
                           => n2576);
   U5991 : MUX2_X1 port map( A => REGISTERS_30_55_port, B => n5819, S => n31, Z
                           => n2575);
   U5992 : MUX2_X1 port map( A => REGISTERS_30_54_port, B => n5820, S => n31, Z
                           => n2574);
   U5993 : MUX2_X1 port map( A => REGISTERS_30_53_port, B => n5821, S => n31, Z
                           => n2573);
   U5994 : MUX2_X1 port map( A => REGISTERS_30_52_port, B => n5822, S => n31, Z
                           => n2572);
   U5995 : MUX2_X1 port map( A => REGISTERS_30_51_port, B => n5823, S => n31, Z
                           => n2571);
   U5996 : MUX2_X1 port map( A => REGISTERS_30_50_port, B => n5824, S => n31, Z
                           => n2570);
   U5997 : MUX2_X1 port map( A => REGISTERS_30_49_port, B => n5825, S => n31, Z
                           => n2569);
   U5998 : MUX2_X1 port map( A => REGISTERS_30_48_port, B => n5826, S => n31, Z
                           => n2568);
   U5999 : MUX2_X1 port map( A => REGISTERS_30_47_port, B => n5827, S => n31, Z
                           => n2567);
   U6000 : MUX2_X1 port map( A => REGISTERS_30_46_port, B => n5828, S => n31, Z
                           => n2566);
   U6001 : MUX2_X1 port map( A => REGISTERS_30_45_port, B => n5829, S => n31, Z
                           => n2565);
   U6002 : MUX2_X1 port map( A => REGISTERS_30_44_port, B => n5830, S => n31, Z
                           => n2564);
   U6003 : MUX2_X1 port map( A => REGISTERS_30_43_port, B => n5831, S => n31, Z
                           => n2563);
   U6004 : MUX2_X1 port map( A => REGISTERS_30_42_port, B => n5832, S => n31, Z
                           => n2562);
   U6005 : MUX2_X1 port map( A => REGISTERS_30_41_port, B => n5833, S => n31, Z
                           => n2561);
   U6006 : MUX2_X1 port map( A => REGISTERS_30_40_port, B => n5834, S => n31, Z
                           => n2560);
   U6007 : MUX2_X1 port map( A => REGISTERS_30_39_port, B => n5835, S => n31, Z
                           => n2559);
   U6008 : MUX2_X1 port map( A => REGISTERS_30_38_port, B => n5836, S => n31, Z
                           => n2558);
   U6009 : MUX2_X1 port map( A => REGISTERS_30_37_port, B => n5837, S => n31, Z
                           => n2557);
   U6010 : MUX2_X1 port map( A => REGISTERS_30_36_port, B => n5838, S => n31, Z
                           => n2556);
   U6011 : MUX2_X1 port map( A => REGISTERS_30_35_port, B => n5839, S => n31, Z
                           => n2555);
   U6012 : MUX2_X1 port map( A => REGISTERS_30_34_port, B => n5840, S => n31, Z
                           => n2554);
   U6013 : MUX2_X1 port map( A => REGISTERS_30_33_port, B => n5841, S => n31, Z
                           => n2553);
   U6014 : MUX2_X1 port map( A => REGISTERS_30_32_port, B => n5842, S => n31, Z
                           => n2552);
   U6015 : MUX2_X1 port map( A => REGISTERS_30_31_port, B => n5843, S => n31, Z
                           => n2551);
   U6016 : MUX2_X1 port map( A => REGISTERS_30_30_port, B => n5844, S => n31, Z
                           => n2550);
   U6017 : MUX2_X1 port map( A => REGISTERS_30_29_port, B => n5845, S => n31, Z
                           => n2549);
   U6018 : MUX2_X1 port map( A => REGISTERS_30_28_port, B => n5846, S => n31, Z
                           => n2548);
   U6019 : MUX2_X1 port map( A => REGISTERS_30_27_port, B => n5847, S => n31, Z
                           => n2547);
   U6020 : MUX2_X1 port map( A => REGISTERS_30_26_port, B => n5848, S => n31, Z
                           => n2546);
   U6021 : MUX2_X1 port map( A => REGISTERS_30_25_port, B => n5849, S => n31, Z
                           => n2545);
   U6022 : MUX2_X1 port map( A => REGISTERS_30_24_port, B => n5850, S => n31, Z
                           => n2544);
   U6023 : MUX2_X1 port map( A => REGISTERS_30_23_port, B => n5851, S => n31, Z
                           => n2543);
   U6024 : MUX2_X1 port map( A => REGISTERS_30_22_port, B => n5852, S => n31, Z
                           => n2542);
   U6025 : MUX2_X1 port map( A => REGISTERS_30_21_port, B => n5853, S => n31, Z
                           => n2541);
   U6026 : MUX2_X1 port map( A => REGISTERS_30_20_port, B => n5854, S => n31, Z
                           => n2540);
   U6027 : MUX2_X1 port map( A => REGISTERS_30_19_port, B => n5855, S => n31, Z
                           => n2539);
   U6028 : MUX2_X1 port map( A => REGISTERS_30_18_port, B => n5856, S => n31, Z
                           => n2538);
   U6029 : MUX2_X1 port map( A => REGISTERS_30_17_port, B => n5857, S => n31, Z
                           => n2537);
   U6030 : MUX2_X1 port map( A => REGISTERS_30_16_port, B => n5858, S => n31, Z
                           => n2536);
   U6031 : MUX2_X1 port map( A => REGISTERS_30_15_port, B => n5859, S => n31, Z
                           => n2535);
   U6032 : MUX2_X1 port map( A => REGISTERS_30_14_port, B => n5860, S => n31, Z
                           => n2534);
   U6033 : MUX2_X1 port map( A => REGISTERS_30_13_port, B => n5861, S => n31, Z
                           => n2533);
   U6034 : MUX2_X1 port map( A => REGISTERS_30_12_port, B => n5862, S => n31, Z
                           => n2532);
   U6035 : MUX2_X1 port map( A => REGISTERS_30_11_port, B => n5863, S => n31, Z
                           => n2531);
   U6036 : MUX2_X1 port map( A => REGISTERS_30_10_port, B => n5864, S => n31, Z
                           => n2530);
   U6037 : MUX2_X1 port map( A => REGISTERS_30_9_port, B => n5865, S => n31, Z 
                           => n2529);
   U6038 : MUX2_X1 port map( A => REGISTERS_30_8_port, B => n5866, S => n31, Z 
                           => n2528);
   U6039 : MUX2_X1 port map( A => REGISTERS_30_7_port, B => n5867, S => n31, Z 
                           => n2527);
   U6040 : MUX2_X1 port map( A => REGISTERS_30_6_port, B => n5868, S => n31, Z 
                           => n2526);
   U6041 : MUX2_X1 port map( A => REGISTERS_30_5_port, B => n5869, S => n31, Z 
                           => n2525);
   U6042 : MUX2_X1 port map( A => REGISTERS_30_4_port, B => n5870, S => n31, Z 
                           => n2524);
   U6043 : MUX2_X1 port map( A => REGISTERS_30_3_port, B => n5871, S => n31, Z 
                           => n2523);
   U6044 : MUX2_X1 port map( A => REGISTERS_30_2_port, B => n5872, S => n31, Z 
                           => n2522);
   U6045 : MUX2_X1 port map( A => REGISTERS_30_1_port, B => n5873, S => n31, Z 
                           => n2521);
   U6046 : MUX2_X1 port map( A => REGISTERS_30_0_port, B => n5874, S => n31, Z 
                           => n2520);
   U6047 : OAI21_X1 port map( B1 => n5888, B2 => n5913, A => n5744, ZN => n5922
                           );
   U6048 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n5916, A3 => ADD_WR(2), ZN
                           => n5888);
   U6049 : INV_X1 port map( A => ADD_WR(0), ZN => n5916);
   U6050 : MUX2_X1 port map( A => REGISTERS_31_63_port, B => n5810, S => n26, Z
                           => n2519);
   U6051 : AND2_X1 port map( A1 => DATAIN(63), A2 => n5744, ZN => n5810);
   U6052 : MUX2_X1 port map( A => REGISTERS_31_62_port, B => n5812, S => n26, Z
                           => n2518);
   U6053 : AND2_X1 port map( A1 => DATAIN(62), A2 => n5744, ZN => n5812);
   U6054 : MUX2_X1 port map( A => REGISTERS_31_61_port, B => n5813, S => n26, Z
                           => n2517);
   U6055 : AND2_X1 port map( A1 => DATAIN(61), A2 => n5744, ZN => n5813);
   U6056 : MUX2_X1 port map( A => REGISTERS_31_60_port, B => n5814, S => n26, Z
                           => n2516);
   U6057 : AND2_X1 port map( A1 => DATAIN(60), A2 => n5744, ZN => n5814);
   U6058 : MUX2_X1 port map( A => REGISTERS_31_59_port, B => n5815, S => n26, Z
                           => n2515);
   U6059 : AND2_X1 port map( A1 => DATAIN(59), A2 => n5744, ZN => n5815);
   U6060 : MUX2_X1 port map( A => REGISTERS_31_58_port, B => n5816, S => n26, Z
                           => n2514);
   U6061 : AND2_X1 port map( A1 => DATAIN(58), A2 => n5744, ZN => n5816);
   U6062 : MUX2_X1 port map( A => REGISTERS_31_57_port, B => n5817, S => n26, Z
                           => n2513);
   U6063 : AND2_X1 port map( A1 => DATAIN(57), A2 => n5744, ZN => n5817);
   U6064 : MUX2_X1 port map( A => REGISTERS_31_56_port, B => n5818, S => n26, Z
                           => n2512);
   U6065 : AND2_X1 port map( A1 => DATAIN(56), A2 => n5744, ZN => n5818);
   U6066 : MUX2_X1 port map( A => REGISTERS_31_55_port, B => n5819, S => n26, Z
                           => n2511);
   U6067 : AND2_X1 port map( A1 => DATAIN(55), A2 => n5744, ZN => n5819);
   U6068 : MUX2_X1 port map( A => REGISTERS_31_54_port, B => n5820, S => n26, Z
                           => n2510);
   U6069 : AND2_X1 port map( A1 => DATAIN(54), A2 => n5744, ZN => n5820);
   U6070 : MUX2_X1 port map( A => REGISTERS_31_53_port, B => n5821, S => n26, Z
                           => n2509);
   U6071 : AND2_X1 port map( A1 => DATAIN(53), A2 => n5744, ZN => n5821);
   U6072 : MUX2_X1 port map( A => REGISTERS_31_52_port, B => n5822, S => n26, Z
                           => n2508);
   U6073 : AND2_X1 port map( A1 => DATAIN(52), A2 => n5744, ZN => n5822);
   U6074 : MUX2_X1 port map( A => REGISTERS_31_51_port, B => n5823, S => n26, Z
                           => n2507);
   U6075 : AND2_X1 port map( A1 => DATAIN(51), A2 => n5744, ZN => n5823);
   U6076 : MUX2_X1 port map( A => REGISTERS_31_50_port, B => n5824, S => n26, Z
                           => n2506);
   U6077 : AND2_X1 port map( A1 => DATAIN(50), A2 => n5744, ZN => n5824);
   U6078 : MUX2_X1 port map( A => REGISTERS_31_49_port, B => n5825, S => n26, Z
                           => n2505);
   U6079 : AND2_X1 port map( A1 => DATAIN(49), A2 => n5744, ZN => n5825);
   U6080 : MUX2_X1 port map( A => REGISTERS_31_48_port, B => n5826, S => n26, Z
                           => n2504);
   U6081 : AND2_X1 port map( A1 => DATAIN(48), A2 => n5744, ZN => n5826);
   U6082 : MUX2_X1 port map( A => REGISTERS_31_47_port, B => n5827, S => n26, Z
                           => n2503);
   U6083 : AND2_X1 port map( A1 => DATAIN(47), A2 => n5744, ZN => n5827);
   U6084 : MUX2_X1 port map( A => REGISTERS_31_46_port, B => n5828, S => n26, Z
                           => n2502);
   U6085 : AND2_X1 port map( A1 => DATAIN(46), A2 => n5744, ZN => n5828);
   U6086 : MUX2_X1 port map( A => REGISTERS_31_45_port, B => n5829, S => n26, Z
                           => n2501);
   U6087 : AND2_X1 port map( A1 => DATAIN(45), A2 => n5744, ZN => n5829);
   U6088 : MUX2_X1 port map( A => REGISTERS_31_44_port, B => n5830, S => n26, Z
                           => n2500);
   U6089 : AND2_X1 port map( A1 => DATAIN(44), A2 => n5744, ZN => n5830);
   U6090 : MUX2_X1 port map( A => REGISTERS_31_43_port, B => n5831, S => n26, Z
                           => n2499);
   U6091 : AND2_X1 port map( A1 => DATAIN(43), A2 => n5744, ZN => n5831);
   U6092 : MUX2_X1 port map( A => REGISTERS_31_42_port, B => n5832, S => n26, Z
                           => n2498);
   U6093 : AND2_X1 port map( A1 => DATAIN(42), A2 => n5744, ZN => n5832);
   U6094 : MUX2_X1 port map( A => REGISTERS_31_41_port, B => n5833, S => n26, Z
                           => n2497);
   U6095 : AND2_X1 port map( A1 => DATAIN(41), A2 => n5744, ZN => n5833);
   U6096 : MUX2_X1 port map( A => REGISTERS_31_40_port, B => n5834, S => n26, Z
                           => n2496);
   U6097 : AND2_X1 port map( A1 => DATAIN(40), A2 => n5744, ZN => n5834);
   U6098 : MUX2_X1 port map( A => REGISTERS_31_39_port, B => n5835, S => n26, Z
                           => n2495);
   U6099 : AND2_X1 port map( A1 => DATAIN(39), A2 => n5744, ZN => n5835);
   U6100 : MUX2_X1 port map( A => REGISTERS_31_38_port, B => n5836, S => n26, Z
                           => n2494);
   U6101 : AND2_X1 port map( A1 => DATAIN(38), A2 => n5744, ZN => n5836);
   U6102 : MUX2_X1 port map( A => REGISTERS_31_37_port, B => n5837, S => n26, Z
                           => n2493);
   U6103 : AND2_X1 port map( A1 => DATAIN(37), A2 => n5744, ZN => n5837);
   U6104 : MUX2_X1 port map( A => REGISTERS_31_36_port, B => n5838, S => n26, Z
                           => n2492);
   U6105 : AND2_X1 port map( A1 => DATAIN(36), A2 => n5744, ZN => n5838);
   U6106 : MUX2_X1 port map( A => REGISTERS_31_35_port, B => n5839, S => n26, Z
                           => n2491);
   U6107 : AND2_X1 port map( A1 => DATAIN(35), A2 => n5744, ZN => n5839);
   U6108 : MUX2_X1 port map( A => REGISTERS_31_34_port, B => n5840, S => n26, Z
                           => n2490);
   U6109 : AND2_X1 port map( A1 => DATAIN(34), A2 => n5744, ZN => n5840);
   U6110 : MUX2_X1 port map( A => REGISTERS_31_33_port, B => n5841, S => n26, Z
                           => n2489);
   U6111 : AND2_X1 port map( A1 => DATAIN(33), A2 => n5744, ZN => n5841);
   U6112 : MUX2_X1 port map( A => REGISTERS_31_32_port, B => n5842, S => n26, Z
                           => n2488);
   U6113 : AND2_X1 port map( A1 => DATAIN(32), A2 => n5744, ZN => n5842);
   U6114 : MUX2_X1 port map( A => REGISTERS_31_31_port, B => n5843, S => n26, Z
                           => n2487);
   U6115 : AND2_X1 port map( A1 => DATAIN(31), A2 => n5744, ZN => n5843);
   U6116 : MUX2_X1 port map( A => REGISTERS_31_30_port, B => n5844, S => n26, Z
                           => n2486);
   U6117 : AND2_X1 port map( A1 => DATAIN(30), A2 => n5744, ZN => n5844);
   U6118 : MUX2_X1 port map( A => REGISTERS_31_29_port, B => n5845, S => n26, Z
                           => n2485);
   U6119 : AND2_X1 port map( A1 => DATAIN(29), A2 => n5744, ZN => n5845);
   U6120 : MUX2_X1 port map( A => REGISTERS_31_28_port, B => n5846, S => n26, Z
                           => n2484);
   U6121 : AND2_X1 port map( A1 => DATAIN(28), A2 => n5744, ZN => n5846);
   U6122 : MUX2_X1 port map( A => REGISTERS_31_27_port, B => n5847, S => n26, Z
                           => n2483);
   U6123 : AND2_X1 port map( A1 => DATAIN(27), A2 => n5744, ZN => n5847);
   U6124 : MUX2_X1 port map( A => REGISTERS_31_26_port, B => n5848, S => n26, Z
                           => n2482);
   U6125 : AND2_X1 port map( A1 => DATAIN(26), A2 => n5744, ZN => n5848);
   U6126 : MUX2_X1 port map( A => REGISTERS_31_25_port, B => n5849, S => n26, Z
                           => n2481);
   U6127 : AND2_X1 port map( A1 => DATAIN(25), A2 => n5744, ZN => n5849);
   U6128 : MUX2_X1 port map( A => REGISTERS_31_24_port, B => n5850, S => n26, Z
                           => n2480);
   U6129 : AND2_X1 port map( A1 => DATAIN(24), A2 => n5744, ZN => n5850);
   U6130 : MUX2_X1 port map( A => REGISTERS_31_23_port, B => n5851, S => n26, Z
                           => n2479);
   U6131 : AND2_X1 port map( A1 => DATAIN(23), A2 => n5744, ZN => n5851);
   U6132 : MUX2_X1 port map( A => REGISTERS_31_22_port, B => n5852, S => n26, Z
                           => n2478);
   U6133 : AND2_X1 port map( A1 => DATAIN(22), A2 => n5744, ZN => n5852);
   U6134 : MUX2_X1 port map( A => REGISTERS_31_21_port, B => n5853, S => n26, Z
                           => n2477);
   U6135 : AND2_X1 port map( A1 => DATAIN(21), A2 => n5744, ZN => n5853);
   U6136 : MUX2_X1 port map( A => REGISTERS_31_20_port, B => n5854, S => n26, Z
                           => n2476);
   U6137 : AND2_X1 port map( A1 => DATAIN(20), A2 => n5744, ZN => n5854);
   U6138 : MUX2_X1 port map( A => REGISTERS_31_19_port, B => n5855, S => n26, Z
                           => n2475);
   U6139 : AND2_X1 port map( A1 => DATAIN(19), A2 => n5744, ZN => n5855);
   U6140 : MUX2_X1 port map( A => REGISTERS_31_18_port, B => n5856, S => n26, Z
                           => n2474);
   U6141 : AND2_X1 port map( A1 => DATAIN(18), A2 => n5744, ZN => n5856);
   U6142 : MUX2_X1 port map( A => REGISTERS_31_17_port, B => n5857, S => n26, Z
                           => n2473);
   U6143 : AND2_X1 port map( A1 => DATAIN(17), A2 => n5744, ZN => n5857);
   U6144 : MUX2_X1 port map( A => REGISTERS_31_16_port, B => n5858, S => n26, Z
                           => n2472);
   U6145 : AND2_X1 port map( A1 => DATAIN(16), A2 => n5744, ZN => n5858);
   U6146 : MUX2_X1 port map( A => REGISTERS_31_15_port, B => n5859, S => n26, Z
                           => n2471);
   U6147 : AND2_X1 port map( A1 => DATAIN(15), A2 => n5744, ZN => n5859);
   U6148 : MUX2_X1 port map( A => REGISTERS_31_14_port, B => n5860, S => n26, Z
                           => n2470);
   U6149 : AND2_X1 port map( A1 => DATAIN(14), A2 => n5744, ZN => n5860);
   U6150 : MUX2_X1 port map( A => REGISTERS_31_13_port, B => n5861, S => n26, Z
                           => n2469);
   U6151 : AND2_X1 port map( A1 => DATAIN(13), A2 => n5744, ZN => n5861);
   U6152 : MUX2_X1 port map( A => REGISTERS_31_12_port, B => n5862, S => n26, Z
                           => n2468);
   U6153 : AND2_X1 port map( A1 => DATAIN(12), A2 => n5744, ZN => n5862);
   U6154 : MUX2_X1 port map( A => REGISTERS_31_11_port, B => n5863, S => n26, Z
                           => n2467);
   U6155 : AND2_X1 port map( A1 => DATAIN(11), A2 => n5744, ZN => n5863);
   U6156 : MUX2_X1 port map( A => REGISTERS_31_10_port, B => n5864, S => n26, Z
                           => n2466);
   U6157 : AND2_X1 port map( A1 => DATAIN(10), A2 => n5744, ZN => n5864);
   U6158 : MUX2_X1 port map( A => REGISTERS_31_9_port, B => n5865, S => n26, Z 
                           => n2465);
   U6159 : AND2_X1 port map( A1 => DATAIN(9), A2 => n5744, ZN => n5865);
   U6160 : MUX2_X1 port map( A => REGISTERS_31_8_port, B => n5866, S => n26, Z 
                           => n2464);
   U6161 : AND2_X1 port map( A1 => DATAIN(8), A2 => n5744, ZN => n5866);
   U6162 : MUX2_X1 port map( A => REGISTERS_31_7_port, B => n5867, S => n26, Z 
                           => n2463);
   U6163 : AND2_X1 port map( A1 => DATAIN(7), A2 => n5744, ZN => n5867);
   U6164 : MUX2_X1 port map( A => REGISTERS_31_6_port, B => n5868, S => n26, Z 
                           => n2462);
   U6165 : AND2_X1 port map( A1 => DATAIN(6), A2 => n5744, ZN => n5868);
   U6166 : MUX2_X1 port map( A => REGISTERS_31_5_port, B => n5869, S => n26, Z 
                           => n2461);
   U6167 : AND2_X1 port map( A1 => DATAIN(5), A2 => n5744, ZN => n5869);
   U6168 : MUX2_X1 port map( A => REGISTERS_31_4_port, B => n5870, S => n26, Z 
                           => n2460);
   U6169 : AND2_X1 port map( A1 => DATAIN(4), A2 => n5744, ZN => n5870);
   U6170 : MUX2_X1 port map( A => REGISTERS_31_3_port, B => n5871, S => n26, Z 
                           => n2459);
   U6171 : AND2_X1 port map( A1 => DATAIN(3), A2 => n5744, ZN => n5871);
   U6172 : MUX2_X1 port map( A => REGISTERS_31_2_port, B => n5872, S => n26, Z 
                           => n2458);
   U6173 : AND2_X1 port map( A1 => DATAIN(2), A2 => n5744, ZN => n5872);
   U6174 : MUX2_X1 port map( A => REGISTERS_31_1_port, B => n5873, S => n26, Z 
                           => n2457);
   U6175 : AND2_X1 port map( A1 => DATAIN(1), A2 => n5744, ZN => n5873);
   U6176 : MUX2_X1 port map( A => REGISTERS_31_0_port, B => n5874, S => n26, Z 
                           => n2456);
   U6177 : OAI21_X1 port map( B1 => n5890, B2 => n5913, A => n5744, ZN => n5923
                           );
   U6178 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n5893, A3 => ADD_WR(4), ZN
                           => n5913);
   U6179 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n5893);
   U6180 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n5890);
   U6181 : AND2_X1 port map( A1 => DATAIN(0), A2 => n5744, ZN => n5874);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Logix_control_rf.all;

entity Logix_control_rf is

   port( rest, enable, clock, call, ret, memory_response, RD1, RD2, WR : in 
         std_logic;  data_in : in std_logic_vector (63 downto 0);  memory_bus :
         inout std_logic_vector (63 downto 0);  address_r_1, address_r_2, 
         address_w : in std_logic_vector (4 downto 0);  out_1, out_2 : out 
         std_logic_vector (63 downto 0);  fill, spill : out std_logic;  addr_1,
         addr_2, addr_r : out std_logic_vector (4 downto 0);  cwp_o : out 
         std_logic_vector (1 downto 0));

end Logix_control_rf;

architecture SYN_Behavioral of Logix_control_rf is

   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X8
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component Logix_control_rf_DW01_incdec_1_DW01_incdec_2
      port( A : in std_logic_vector (31 downto 0);  INC_DEC : in std_logic;  
            SUM : out std_logic_vector (31 downto 0));
   end component;
   
   component Logix_control_rf_DW01_incdec_0_DW01_incdec_1
      port( A : in std_logic_vector (31 downto 0);  INC_DEC : in std_logic;  
            SUM : out std_logic_vector (31 downto 0));
   end component;
   
   component register_file_address_length5_Data_parallelism64
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal fill_port, spill_port, addr_1_4_port, addr_1_3_port, addr_1_2_port, 
      addr_1_1_port, addr_2_4_port, addr_2_3_port, addr_2_2_port, addr_2_1_port
      , addr_r_4_port, addr_r_3_port, addr_r_2_port, addr_r_1_port, 
      cwp_o_1_port, rest_s, cansave_31_port, cansave_30_port, cansave_29_port, 
      cansave_28_port, cansave_27_port, cansave_26_port, cansave_25_port, 
      cansave_24_port, cansave_23_port, cansave_22_port, cansave_21_port, 
      cansave_20_port, cansave_19_port, cansave_18_port, cansave_17_port, 
      cansave_16_port, cansave_15_port, cansave_14_port, cansave_13_port, 
      cansave_12_port, cansave_11_port, cansave_10_port, cansave_9_port, 
      cansave_8_port, cansave_7_port, cansave_6_port, cansave_5_port, 
      cansave_4_port, cansave_3_port, cansave_2_port, cansave_1_port, 
      cansave_0_port, canrestore_31_port, canrestore_30_port, 
      canrestore_29_port, canrestore_28_port, canrestore_27_port, 
      canrestore_26_port, canrestore_25_port, canrestore_24_port, 
      canrestore_23_port, canrestore_22_port, canrestore_21_port, 
      canrestore_20_port, canrestore_19_port, canrestore_18_port, 
      canrestore_17_port, canrestore_16_port, canrestore_15_port, 
      canrestore_14_port, canrestore_13_port, canrestore_12_port, 
      canrestore_11_port, canrestore_10_port, canrestore_9_port, 
      canrestore_8_port, canrestore_7_port, canrestore_6_port, 
      canrestore_5_port, canrestore_4_port, canrestore_3_port, 
      canrestore_2_port, canrestore_1_port, canrestore_0_port, N246, N247, N248
      , N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
      N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, 
      N273, N274, N275, N276, N277, N645, N646, N647, N648, N649, N650, N651, 
      N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, 
      N664, N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675, 
      N676, N1006, N1274, U3_U6_Z_0, n273_port, n402, n403, n404, n405, n406, 
      n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, 
      n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
      n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, 
      n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, 
      n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, 
      n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, 
      n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, 
      n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, 
      n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, 
      n645_port, n646_port, n647_port, n648_port, n649_port, n650_port, 
      n651_port, n652_port, n653_port, n654_port, n655_port, n656_port, 
      n657_port, n658_port, n659_port, n660_port, n661_port, n662_port, 
      n663_port, n664_port, n665_port, n666_port, n667_port, n668_port, 
      n669_port, n670_port, n671_port, n672_port, n673_port, n674_port, 
      n675_port, n676_port, n677, n678, n679, n680, n681, n682, n683, n684, 
      n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, 
      n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, 
      n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, 
      n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, 
      n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, 
      n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, 
      n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, 
      n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
      n793, n794, n795, r339_LEQ, n799, n800, n801, n802, n803, n804, n805, 
      n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, 
      n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, 
      n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, 
      n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, 
      n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, 
      n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, 
      n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, 
      n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, 
      n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, 
      n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, 
      n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, 
      n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, 
      n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, 
      n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, 
      n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, 
      n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, 
      n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006_port, n1007, 
      n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
      n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
      n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, 
      n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, 
      n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, 
      n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, 
      n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, 
      n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, 
      n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, 
      n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, 
      n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, 
      n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, 
      n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, 
      n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, 
      n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, 
      n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, 
      n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, 
      n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, 
      n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, 
      n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, 
      n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, 
      n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
      n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, 
      n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, 
      n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, 
      n1258, n1259, n1260, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, 
      n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3066, 
      n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, 
      n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, n_3083, n_3084, 
      n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091, n_3092, n_3093, 
      n_3094, n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, 
      n_3103, n_3104, n_3105, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, 
      n_3112, n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120 : 
      std_logic;

begin
   fill <= fill_port;
   spill <= spill_port;
   addr_1 <= ( addr_1_4_port, addr_1_3_port, addr_1_2_port, addr_1_1_port, 
      address_r_1(0) );
   addr_2 <= ( addr_2_4_port, addr_2_3_port, addr_2_2_port, addr_2_1_port, 
      address_r_2(0) );
   addr_r <= ( addr_r_4_port, addr_r_3_port, addr_r_2_port, addr_r_1_port, 
      address_w(0) );
   cwp_o <= ( cwp_o_1_port, N1274 );
   
   next_state_reg_0_inst : DFF_X1 port map( D => n794, CK => n869, Q => n_3052,
                           QN => n1131);
   cansave_reg_0_inst : DFF_X1 port map( D => n795, CK => n868, Q => 
                           cansave_0_port, QN => n466);
   next_state_reg_1_inst : DFF_X1 port map( D => n794, CK => n869, Q => n_3053,
                           QN => n1132);
   rest_s_reg : DFF_X1 port map( D => N1006, CK => n869, Q => rest_s, QN => 
                           n_3054);
   canrestore_reg_0_inst : DFF_X1 port map( D => n793, CK => n868, Q => 
                           canrestore_0_port, QN => n465);
   canrestore_reg_31_inst : DFF_X1 port map( D => n792, CK => n868, Q => 
                           canrestore_31_port, QN => n464);
   canrestore_reg_30_inst : DFF_X1 port map( D => n791, CK => n868, Q => 
                           canrestore_30_port, QN => n463);
   canrestore_reg_29_inst : DFF_X1 port map( D => n790, CK => n868, Q => 
                           canrestore_29_port, QN => n462);
   canrestore_reg_28_inst : DFF_X1 port map( D => n789, CK => n868, Q => 
                           canrestore_28_port, QN => n461);
   canrestore_reg_27_inst : DFF_X1 port map( D => n788, CK => n868, Q => 
                           canrestore_27_port, QN => n460);
   canrestore_reg_26_inst : DFF_X1 port map( D => n787, CK => n868, Q => 
                           canrestore_26_port, QN => n459);
   canrestore_reg_25_inst : DFF_X1 port map( D => n786, CK => n868, Q => 
                           canrestore_25_port, QN => n458);
   canrestore_reg_24_inst : DFF_X1 port map( D => n785, CK => n868, Q => 
                           canrestore_24_port, QN => n457);
   canrestore_reg_23_inst : DFF_X1 port map( D => n784, CK => n868, Q => 
                           canrestore_23_port, QN => n456);
   canrestore_reg_22_inst : DFF_X1 port map( D => n783, CK => n868, Q => 
                           canrestore_22_port, QN => n455);
   canrestore_reg_21_inst : DFF_X1 port map( D => n782, CK => n868, Q => 
                           canrestore_21_port, QN => n454);
   canrestore_reg_20_inst : DFF_X1 port map( D => n781, CK => n868, Q => 
                           canrestore_20_port, QN => n453);
   canrestore_reg_19_inst : DFF_X1 port map( D => n780, CK => n868, Q => 
                           canrestore_19_port, QN => n452);
   canrestore_reg_18_inst : DFF_X1 port map( D => n779, CK => n868, Q => 
                           canrestore_18_port, QN => n451);
   canrestore_reg_17_inst : DFF_X1 port map( D => n778, CK => n868, Q => 
                           canrestore_17_port, QN => n450);
   canrestore_reg_16_inst : DFF_X1 port map( D => n777, CK => n868, Q => 
                           canrestore_16_port, QN => n449);
   canrestore_reg_15_inst : DFF_X1 port map( D => n776, CK => n868, Q => 
                           canrestore_15_port, QN => n448);
   canrestore_reg_14_inst : DFF_X1 port map( D => n775, CK => n868, Q => 
                           canrestore_14_port, QN => n447);
   canrestore_reg_13_inst : DFF_X1 port map( D => n774, CK => n868, Q => 
                           canrestore_13_port, QN => n446);
   canrestore_reg_12_inst : DFF_X1 port map( D => n773, CK => n868, Q => 
                           canrestore_12_port, QN => n445);
   canrestore_reg_11_inst : DFF_X1 port map( D => n772, CK => n868, Q => 
                           canrestore_11_port, QN => n444);
   canrestore_reg_10_inst : DFF_X1 port map( D => n771, CK => n868, Q => 
                           canrestore_10_port, QN => n443);
   canrestore_reg_9_inst : DFF_X1 port map( D => n770, CK => n868, Q => 
                           canrestore_9_port, QN => n442);
   canrestore_reg_8_inst : DFF_X1 port map( D => n769, CK => n868, Q => 
                           canrestore_8_port, QN => n441);
   canrestore_reg_7_inst : DFF_X1 port map( D => n768, CK => n868, Q => 
                           canrestore_7_port, QN => n440);
   canrestore_reg_6_inst : DFF_X1 port map( D => n767, CK => n868, Q => 
                           canrestore_6_port, QN => n439);
   canrestore_reg_5_inst : DFF_X1 port map( D => n766, CK => n868, Q => 
                           canrestore_5_port, QN => n438);
   canrestore_reg_4_inst : DFF_X1 port map( D => n765, CK => n868, Q => 
                           canrestore_4_port, QN => n437);
   canrestore_reg_3_inst : DFF_X1 port map( D => n764, CK => n868, Q => 
                           canrestore_3_port, QN => n436);
   canrestore_reg_2_inst : DFF_X1 port map( D => n763, CK => n868, Q => 
                           canrestore_2_port, QN => n435);
   canrestore_reg_1_inst : DFF_X1 port map( D => n762, CK => n868, Q => 
                           canrestore_1_port, QN => n434);
   cwp_reg_0_inst : DFF_X1 port map( D => n761, CK => n868, Q => N1274, QN => 
                           n433);
   cansave_reg_1_inst : DFF_X1 port map( D => n760, CK => n868, Q => 
                           cansave_1_port, QN => n432);
   cansave_reg_31_inst : DFF_X1 port map( D => n759, CK => n868, Q => 
                           cansave_31_port, QN => n431);
   cansave_reg_2_inst : DFF_X1 port map( D => n758, CK => n868, Q => 
                           cansave_2_port, QN => n430);
   cansave_reg_30_inst : DFF_X1 port map( D => n757, CK => n868, Q => 
                           cansave_30_port, QN => n429);
   cansave_reg_29_inst : DFF_X1 port map( D => n756, CK => n868, Q => 
                           cansave_29_port, QN => n428);
   cansave_reg_28_inst : DFF_X1 port map( D => n755, CK => n868, Q => 
                           cansave_28_port, QN => n427);
   cansave_reg_27_inst : DFF_X1 port map( D => n754, CK => n868, Q => 
                           cansave_27_port, QN => n426);
   cansave_reg_26_inst : DFF_X1 port map( D => n753, CK => n868, Q => 
                           cansave_26_port, QN => n425);
   cansave_reg_25_inst : DFF_X1 port map( D => n752, CK => n868, Q => 
                           cansave_25_port, QN => n424);
   cansave_reg_24_inst : DFF_X1 port map( D => n751, CK => n868, Q => 
                           cansave_24_port, QN => n423);
   cansave_reg_23_inst : DFF_X1 port map( D => n750, CK => n868, Q => 
                           cansave_23_port, QN => n422);
   cansave_reg_22_inst : DFF_X1 port map( D => n749, CK => n868, Q => 
                           cansave_22_port, QN => n421);
   cansave_reg_21_inst : DFF_X1 port map( D => n748, CK => n868, Q => 
                           cansave_21_port, QN => n420);
   cansave_reg_20_inst : DFF_X1 port map( D => n747, CK => n868, Q => 
                           cansave_20_port, QN => n419);
   cansave_reg_19_inst : DFF_X1 port map( D => n746, CK => n868, Q => 
                           cansave_19_port, QN => n418);
   cansave_reg_18_inst : DFF_X1 port map( D => n745, CK => n868, Q => 
                           cansave_18_port, QN => n417);
   cansave_reg_17_inst : DFF_X1 port map( D => n744, CK => n868, Q => 
                           cansave_17_port, QN => n416);
   cansave_reg_16_inst : DFF_X1 port map( D => n743, CK => n868, Q => 
                           cansave_16_port, QN => n415);
   cansave_reg_15_inst : DFF_X1 port map( D => n742, CK => n868, Q => 
                           cansave_15_port, QN => n414);
   cansave_reg_14_inst : DFF_X1 port map( D => n741, CK => n868, Q => 
                           cansave_14_port, QN => n413);
   cansave_reg_13_inst : DFF_X1 port map( D => n740, CK => n868, Q => 
                           cansave_13_port, QN => n412);
   cansave_reg_12_inst : DFF_X1 port map( D => n739, CK => n868, Q => 
                           cansave_12_port, QN => n411);
   cansave_reg_11_inst : DFF_X1 port map( D => n738, CK => n868, Q => 
                           cansave_11_port, QN => n410);
   cansave_reg_10_inst : DFF_X1 port map( D => n737, CK => n868, Q => 
                           cansave_10_port, QN => n409);
   cansave_reg_9_inst : DFF_X1 port map( D => n736, CK => n868, Q => 
                           cansave_9_port, QN => n408);
   cansave_reg_8_inst : DFF_X1 port map( D => n735, CK => n868, Q => 
                           cansave_8_port, QN => n407);
   cansave_reg_7_inst : DFF_X1 port map( D => n734, CK => n868, Q => 
                           cansave_7_port, QN => n406);
   cansave_reg_6_inst : DFF_X1 port map( D => n733, CK => n868, Q => 
                           cansave_6_port, QN => n405);
   cansave_reg_5_inst : DFF_X1 port map( D => n732, CK => n868, Q => 
                           cansave_5_port, QN => n404);
   cansave_reg_4_inst : DFF_X1 port map( D => n731, CK => n868, Q => 
                           cansave_4_port, QN => n403);
   cansave_reg_3_inst : DFF_X1 port map( D => n730, CK => n868, Q => 
                           cansave_3_port, QN => n402);
   next_state_reg_2_inst : DFF_X1 port map( D => n729, CK => n869, Q => n799, 
                           QN => n1130);
   memory_bus_reg_1_inst : DFF_X1 port map( D => n728, CK => n868, Q => n1133, 
                           QN => n_3055);
   memory_bus_tri_enable_reg_1_inst : DFF_X1 port map( D => n727, CK => n868, Q
                           => n1134, QN => n829);
   memory_bus_reg_14_inst : DFF_X1 port map( D => n726, CK => n868, Q => n1135,
                           QN => n_3056);
   memory_bus_tri_enable_reg_14_inst : DFF_X1 port map( D => n725, CK => n868, 
                           Q => n1136, QN => n830);
   memory_bus_reg_13_inst : DFF_X1 port map( D => n724, CK => n868, Q => n1137,
                           QN => n_3057);
   memory_bus_tri_enable_reg_13_inst : DFF_X1 port map( D => n723, CK => n868, 
                           Q => n1138, QN => n831);
   memory_bus_reg_12_inst : DFF_X1 port map( D => n722, CK => n868, Q => n1139,
                           QN => n_3058);
   memory_bus_tri_enable_reg_12_inst : DFF_X1 port map( D => n721, CK => n868, 
                           Q => n1140, QN => n832);
   memory_bus_reg_11_inst : DFF_X1 port map( D => n720, CK => n868, Q => n1141,
                           QN => n_3059);
   memory_bus_tri_enable_reg_11_inst : DFF_X1 port map( D => n719, CK => n868, 
                           Q => n1142, QN => n833);
   memory_bus_reg_10_inst : DFF_X1 port map( D => n718, CK => n868, Q => n1143,
                           QN => n_3060);
   memory_bus_tri_enable_reg_10_inst : DFF_X1 port map( D => n717, CK => n868, 
                           Q => n1144, QN => n834);
   memory_bus_reg_9_inst : DFF_X1 port map( D => n716, CK => n868, Q => n1145, 
                           QN => n_3061);
   memory_bus_tri_enable_reg_9_inst : DFF_X1 port map( D => n715, CK => n868, Q
                           => n1146, QN => n835);
   memory_bus_reg_8_inst : DFF_X1 port map( D => n714, CK => n868, Q => n1147, 
                           QN => n_3062);
   memory_bus_tri_enable_reg_8_inst : DFF_X1 port map( D => n713, CK => n868, Q
                           => n1148, QN => n836);
   memory_bus_reg_7_inst : DFF_X1 port map( D => n712, CK => n868, Q => n1149, 
                           QN => n_3063);
   memory_bus_tri_enable_reg_7_inst : DFF_X1 port map( D => n711, CK => n868, Q
                           => n1150, QN => n837);
   memory_bus_reg_6_inst : DFF_X1 port map( D => n710, CK => n868, Q => n1151, 
                           QN => n_3064);
   memory_bus_tri_enable_reg_6_inst : DFF_X1 port map( D => n709, CK => n868, Q
                           => n1152, QN => n838);
   memory_bus_reg_5_inst : DFF_X1 port map( D => n708, CK => n868, Q => n1153, 
                           QN => n_3065);
   memory_bus_tri_enable_reg_5_inst : DFF_X1 port map( D => n707, CK => n868, Q
                           => n1154, QN => n839);
   memory_bus_reg_4_inst : DFF_X1 port map( D => n706, CK => n868, Q => n1155, 
                           QN => n_3066);
   memory_bus_tri_enable_reg_4_inst : DFF_X1 port map( D => n705, CK => n868, Q
                           => n1156, QN => n840);
   memory_bus_reg_3_inst : DFF_X1 port map( D => n704, CK => n868, Q => n1157, 
                           QN => n_3067);
   memory_bus_tri_enable_reg_3_inst : DFF_X1 port map( D => n703, CK => n868, Q
                           => n1158, QN => n841);
   memory_bus_reg_2_inst : DFF_X1 port map( D => n702, CK => n868, Q => n1159, 
                           QN => n_3068);
   memory_bus_tri_enable_reg_2_inst : DFF_X1 port map( D => n701, CK => n868, Q
                           => n1160, QN => n842);
   memory_bus_tri_enable_reg_15_inst : DFF_X1 port map( D => n700, CK => n868, 
                           Q => n1161, QN => n843);
   memory_bus_reg_15_inst : DFF_X1 port map( D => n699, CK => n868, Q => n1162,
                           QN => n_3069);
   memory_bus_tri_enable_reg_16_inst : DFF_X1 port map( D => n698, CK => n868, 
                           Q => n1163, QN => n844);
   memory_bus_reg_16_inst : DFF_X1 port map( D => n697, CK => n868, Q => n1164,
                           QN => n_3070);
   memory_bus_tri_enable_reg_17_inst : DFF_X1 port map( D => n696, CK => n868, 
                           Q => n1165, QN => n845);
   memory_bus_reg_17_inst : DFF_X1 port map( D => n695, CK => n868, Q => n1166,
                           QN => n_3071);
   memory_bus_tri_enable_reg_18_inst : DFF_X1 port map( D => n694, CK => n868, 
                           Q => n1167, QN => n846);
   memory_bus_reg_18_inst : DFF_X1 port map( D => n693, CK => n868, Q => n1168,
                           QN => n_3072);
   memory_bus_tri_enable_reg_19_inst : DFF_X1 port map( D => n692, CK => n868, 
                           Q => n1169, QN => n847);
   memory_bus_reg_19_inst : DFF_X1 port map( D => n691, CK => n868, Q => n1170,
                           QN => n_3073);
   memory_bus_tri_enable_reg_20_inst : DFF_X1 port map( D => n690, CK => n868, 
                           Q => n1171, QN => n848);
   memory_bus_reg_20_inst : DFF_X1 port map( D => n689, CK => n868, Q => n1172,
                           QN => n_3074);
   memory_bus_tri_enable_reg_21_inst : DFF_X1 port map( D => n688, CK => n868, 
                           Q => n1173, QN => n849);
   memory_bus_reg_21_inst : DFF_X1 port map( D => n687, CK => n868, Q => n1174,
                           QN => n_3075);
   memory_bus_tri_enable_reg_22_inst : DFF_X1 port map( D => n686, CK => n868, 
                           Q => n1175, QN => n850);
   memory_bus_reg_22_inst : DFF_X1 port map( D => n685, CK => n868, Q => n1176,
                           QN => n_3076);
   memory_bus_tri_enable_reg_23_inst : DFF_X1 port map( D => n684, CK => n868, 
                           Q => n1177, QN => n851);
   memory_bus_reg_23_inst : DFF_X1 port map( D => n683, CK => n868, Q => n1178,
                           QN => n_3077);
   memory_bus_tri_enable_reg_24_inst : DFF_X1 port map( D => n682, CK => n868, 
                           Q => n1179, QN => n852);
   memory_bus_reg_24_inst : DFF_X1 port map( D => n681, CK => n868, Q => n1180,
                           QN => n_3078);
   memory_bus_tri_enable_reg_25_inst : DFF_X1 port map( D => n680, CK => n868, 
                           Q => n1181, QN => n853);
   memory_bus_reg_25_inst : DFF_X1 port map( D => n679, CK => n868, Q => n1182,
                           QN => n_3079);
   memory_bus_tri_enable_reg_26_inst : DFF_X1 port map( D => n678, CK => n868, 
                           Q => n1183, QN => n854);
   memory_bus_reg_26_inst : DFF_X1 port map( D => n677, CK => n868, Q => n1184,
                           QN => n_3080);
   memory_bus_tri_enable_reg_27_inst : DFF_X1 port map( D => n676_port, CK => 
                           n868, Q => n1185, QN => n855);
   memory_bus_reg_27_inst : DFF_X1 port map( D => n675_port, CK => n868, Q => 
                           n1186, QN => n_3081);
   memory_bus_tri_enable_reg_28_inst : DFF_X1 port map( D => n674_port, CK => 
                           n868, Q => n1187, QN => n856);
   memory_bus_reg_28_inst : DFF_X1 port map( D => n673_port, CK => n868, Q => 
                           n1188, QN => n_3082);
   memory_bus_tri_enable_reg_29_inst : DFF_X1 port map( D => n672_port, CK => 
                           n868, Q => n1189, QN => n857);
   memory_bus_reg_29_inst : DFF_X1 port map( D => n671_port, CK => n868, Q => 
                           n1190, QN => n_3083);
   memory_bus_tri_enable_reg_30_inst : DFF_X1 port map( D => n670_port, CK => 
                           n868, Q => n1191, QN => n858);
   memory_bus_reg_30_inst : DFF_X1 port map( D => n669_port, CK => n868, Q => 
                           n1192, QN => n_3084);
   memory_bus_tri_enable_reg_31_inst : DFF_X1 port map( D => n668_port, CK => 
                           n868, Q => n1193, QN => n859);
   memory_bus_reg_31_inst : DFF_X1 port map( D => n667_port, CK => n868, Q => 
                           n1194, QN => n_3085);
   memory_bus_tri_enable_reg_32_inst : DFF_X1 port map( D => n666_port, CK => 
                           n868, Q => n1195, QN => n860);
   memory_bus_reg_32_inst : DFF_X1 port map( D => n665_port, CK => n868, Q => 
                           n1196, QN => n_3086);
   memory_bus_tri_enable_reg_33_inst : DFF_X1 port map( D => n664_port, CK => 
                           n868, Q => n1197, QN => n861);
   memory_bus_reg_33_inst : DFF_X1 port map( D => n663_port, CK => n868, Q => 
                           n1198, QN => n_3087);
   memory_bus_tri_enable_reg_34_inst : DFF_X1 port map( D => n662_port, CK => 
                           n868, Q => n1199, QN => n862);
   memory_bus_reg_34_inst : DFF_X1 port map( D => n661_port, CK => n868, Q => 
                           n1200, QN => n_3088);
   memory_bus_tri_enable_reg_35_inst : DFF_X1 port map( D => n660_port, CK => 
                           n868, Q => n1201, QN => n863);
   memory_bus_reg_35_inst : DFF_X1 port map( D => n659_port, CK => n868, Q => 
                           n1202, QN => n_3089);
   memory_bus_tri_enable_reg_36_inst : DFF_X1 port map( D => n658_port, CK => 
                           n869, Q => n1203, QN => n800);
   memory_bus_reg_36_inst : DFF_X1 port map( D => n657_port, CK => n868, Q => 
                           n1204, QN => n_3090);
   memory_bus_tri_enable_reg_37_inst : DFF_X1 port map( D => n656_port, CK => 
                           n869, Q => n1205, QN => n801);
   memory_bus_reg_37_inst : DFF_X1 port map( D => n655_port, CK => n868, Q => 
                           n1206, QN => n_3091);
   memory_bus_tri_enable_reg_38_inst : DFF_X1 port map( D => n654_port, CK => 
                           n869, Q => n1207, QN => n802);
   memory_bus_reg_38_inst : DFF_X1 port map( D => n653_port, CK => n868, Q => 
                           n1208, QN => n_3092);
   memory_bus_tri_enable_reg_39_inst : DFF_X1 port map( D => n652_port, CK => 
                           n869, Q => n1209, QN => n803);
   memory_bus_reg_39_inst : DFF_X1 port map( D => n651_port, CK => n868, Q => 
                           n1210, QN => n_3093);
   memory_bus_tri_enable_reg_40_inst : DFF_X1 port map( D => n650_port, CK => 
                           n869, Q => n1211, QN => n804);
   memory_bus_reg_40_inst : DFF_X1 port map( D => n649_port, CK => n868, Q => 
                           n1212, QN => n_3094);
   memory_bus_tri_enable_reg_41_inst : DFF_X1 port map( D => n648_port, CK => 
                           n869, Q => n1213, QN => n805);
   memory_bus_reg_41_inst : DFF_X1 port map( D => n647_port, CK => n868, Q => 
                           n1214, QN => n_3095);
   memory_bus_tri_enable_reg_42_inst : DFF_X1 port map( D => n646_port, CK => 
                           n869, Q => n1215, QN => n806);
   memory_bus_reg_42_inst : DFF_X1 port map( D => n645_port, CK => n868, Q => 
                           n1216, QN => n_3096);
   memory_bus_tri_enable_reg_43_inst : DFF_X1 port map( D => n644, CK => n869, 
                           Q => n1217, QN => n807);
   memory_bus_reg_43_inst : DFF_X1 port map( D => n643, CK => n868, Q => n1218,
                           QN => n_3097);
   memory_bus_tri_enable_reg_44_inst : DFF_X1 port map( D => n642, CK => n869, 
                           Q => n1219, QN => n808);
   memory_bus_reg_44_inst : DFF_X1 port map( D => n641, CK => n868, Q => n1220,
                           QN => n_3098);
   memory_bus_tri_enable_reg_45_inst : DFF_X1 port map( D => n640, CK => n869, 
                           Q => n1221, QN => n809);
   memory_bus_reg_45_inst : DFF_X1 port map( D => n639, CK => n868, Q => n1222,
                           QN => n_3099);
   memory_bus_tri_enable_reg_46_inst : DFF_X1 port map( D => n638, CK => n869, 
                           Q => n1223, QN => n810);
   memory_bus_reg_46_inst : DFF_X1 port map( D => n637, CK => n868, Q => n1224,
                           QN => n_3100);
   memory_bus_tri_enable_reg_47_inst : DFF_X1 port map( D => n636, CK => n869, 
                           Q => n1225, QN => n811);
   memory_bus_reg_47_inst : DFF_X1 port map( D => n635, CK => n868, Q => n1226,
                           QN => n_3101);
   memory_bus_tri_enable_reg_48_inst : DFF_X1 port map( D => n634, CK => n869, 
                           Q => n1227, QN => n812);
   memory_bus_reg_48_inst : DFF_X1 port map( D => n633, CK => n868, Q => n1228,
                           QN => n_3102);
   memory_bus_tri_enable_reg_49_inst : DFF_X1 port map( D => n632, CK => n869, 
                           Q => n1229, QN => n813);
   memory_bus_reg_49_inst : DFF_X1 port map( D => n631, CK => n868, Q => n1230,
                           QN => n_3103);
   memory_bus_tri_enable_reg_50_inst : DFF_X1 port map( D => n630, CK => n869, 
                           Q => n1231, QN => n814);
   memory_bus_reg_50_inst : DFF_X1 port map( D => n629, CK => n868, Q => n1232,
                           QN => n_3104);
   memory_bus_tri_enable_reg_51_inst : DFF_X1 port map( D => n628, CK => n869, 
                           Q => n1233, QN => n815);
   memory_bus_reg_51_inst : DFF_X1 port map( D => n627, CK => n868, Q => n1234,
                           QN => n_3105);
   memory_bus_tri_enable_reg_52_inst : DFF_X1 port map( D => n626, CK => n869, 
                           Q => n1235, QN => n816);
   memory_bus_reg_52_inst : DFF_X1 port map( D => n625, CK => n868, Q => n1236,
                           QN => n_3106);
   memory_bus_tri_enable_reg_53_inst : DFF_X1 port map( D => n624, CK => n869, 
                           Q => n1237, QN => n817);
   memory_bus_reg_53_inst : DFF_X1 port map( D => n623, CK => n868, Q => n1238,
                           QN => n_3107);
   memory_bus_tri_enable_reg_54_inst : DFF_X1 port map( D => n622, CK => n869, 
                           Q => n1239, QN => n818);
   memory_bus_reg_54_inst : DFF_X1 port map( D => n621, CK => n868, Q => n1240,
                           QN => n_3108);
   memory_bus_tri_enable_reg_55_inst : DFF_X1 port map( D => n620, CK => n869, 
                           Q => n1241, QN => n819);
   memory_bus_reg_55_inst : DFF_X1 port map( D => n619, CK => n868, Q => n1242,
                           QN => n_3109);
   memory_bus_tri_enable_reg_56_inst : DFF_X1 port map( D => n618, CK => n869, 
                           Q => n1243, QN => n820);
   memory_bus_reg_56_inst : DFF_X1 port map( D => n617, CK => n868, Q => n1244,
                           QN => n_3110);
   memory_bus_tri_enable_reg_57_inst : DFF_X1 port map( D => n616, CK => n869, 
                           Q => n1245, QN => n821);
   memory_bus_reg_57_inst : DFF_X1 port map( D => n615, CK => n868, Q => n1246,
                           QN => n_3111);
   memory_bus_tri_enable_reg_58_inst : DFF_X1 port map( D => n614, CK => n869, 
                           Q => n1247, QN => n822);
   memory_bus_reg_58_inst : DFF_X1 port map( D => n613, CK => n868, Q => n1248,
                           QN => n_3112);
   memory_bus_tri_enable_reg_59_inst : DFF_X1 port map( D => n612, CK => n869, 
                           Q => n1249, QN => n823);
   memory_bus_reg_59_inst : DFF_X1 port map( D => n611, CK => n868, Q => n1250,
                           QN => n_3113);
   memory_bus_tri_enable_reg_60_inst : DFF_X1 port map( D => n610, CK => n869, 
                           Q => n1251, QN => n824);
   memory_bus_reg_60_inst : DFF_X1 port map( D => n609, CK => n868, Q => n1252,
                           QN => n_3114);
   memory_bus_tri_enable_reg_61_inst : DFF_X1 port map( D => n608, CK => n869, 
                           Q => n1253, QN => n825);
   memory_bus_reg_61_inst : DFF_X1 port map( D => n607, CK => n868, Q => n1254,
                           QN => n_3115);
   memory_bus_tri_enable_reg_62_inst : DFF_X1 port map( D => n606, CK => n869, 
                           Q => n1255, QN => n826);
   memory_bus_reg_62_inst : DFF_X1 port map( D => n605, CK => n868, Q => n1256,
                           QN => n_3116);
   memory_bus_tri_enable_reg_63_inst : DFF_X1 port map( D => n604, CK => n869, 
                           Q => n1257, QN => n827);
   memory_bus_reg_63_inst : DFF_X1 port map( D => n603, CK => n868, Q => n1258,
                           QN => n_3117);
   memory_bus_tri_enable_reg_0_inst : DFF_X1 port map( D => n602, CK => n869, Q
                           => n1259, QN => n828);
   memory_bus_reg_0_inst : DFF_X1 port map( D => n601, CK => n868, Q => n1260, 
                           QN => n_3118);
   cwp_reg_1_inst : DFF_X1 port map( D => n600, CK => n868, Q => cwp_o_1_port, 
                           QN => n273_port);
   spill_reg : DFF_X1 port map( D => n599, CK => n868, Q => spill_port, QN => 
                           n_3119);
   fill_reg : DFF_X1 port map( D => n598, CK => n868, Q => fill_port, QN => 
                           n_3120);
   L : register_file_address_length5_Data_parallelism64 port map( CLK => n868, 
                           RESET => rest_s, ENABLE => enable, RD1 => RD1, RD2 
                           => RD2, WR => WR, ADD_WR(4) => addr_r_4_port, 
                           ADD_WR(3) => addr_r_3_port, ADD_WR(2) => 
                           addr_r_2_port, ADD_WR(1) => addr_r_1_port, ADD_WR(0)
                           => address_w(0), ADD_RD1(4) => addr_1_4_port, 
                           ADD_RD1(3) => addr_1_3_port, ADD_RD1(2) => 
                           addr_1_2_port, ADD_RD1(1) => addr_1_1_port, 
                           ADD_RD1(0) => address_r_1(0), ADD_RD2(4) => 
                           addr_2_4_port, ADD_RD2(3) => addr_2_3_port, 
                           ADD_RD2(2) => addr_2_2_port, ADD_RD2(1) => 
                           addr_2_1_port, ADD_RD2(0) => address_r_2(0), 
                           DATAIN(63) => data_in(63), DATAIN(62) => data_in(62)
                           , DATAIN(61) => data_in(61), DATAIN(60) => 
                           data_in(60), DATAIN(59) => data_in(59), DATAIN(58) 
                           => data_in(58), DATAIN(57) => data_in(57), 
                           DATAIN(56) => data_in(56), DATAIN(55) => data_in(55)
                           , DATAIN(54) => data_in(54), DATAIN(53) => 
                           data_in(53), DATAIN(52) => data_in(52), DATAIN(51) 
                           => data_in(51), DATAIN(50) => data_in(50), 
                           DATAIN(49) => data_in(49), DATAIN(48) => data_in(48)
                           , DATAIN(47) => data_in(47), DATAIN(46) => 
                           data_in(46), DATAIN(45) => data_in(45), DATAIN(44) 
                           => data_in(44), DATAIN(43) => data_in(43), 
                           DATAIN(42) => data_in(42), DATAIN(41) => data_in(41)
                           , DATAIN(40) => data_in(40), DATAIN(39) => 
                           data_in(39), DATAIN(38) => data_in(38), DATAIN(37) 
                           => data_in(37), DATAIN(36) => data_in(36), 
                           DATAIN(35) => data_in(35), DATAIN(34) => data_in(34)
                           , DATAIN(33) => data_in(33), DATAIN(32) => 
                           data_in(32), DATAIN(31) => data_in(31), DATAIN(30) 
                           => data_in(30), DATAIN(29) => data_in(29), 
                           DATAIN(28) => data_in(28), DATAIN(27) => data_in(27)
                           , DATAIN(26) => data_in(26), DATAIN(25) => 
                           data_in(25), DATAIN(24) => data_in(24), DATAIN(23) 
                           => data_in(23), DATAIN(22) => data_in(22), 
                           DATAIN(21) => data_in(21), DATAIN(20) => data_in(20)
                           , DATAIN(19) => data_in(19), DATAIN(18) => 
                           data_in(18), DATAIN(17) => data_in(17), DATAIN(16) 
                           => data_in(16), DATAIN(15) => data_in(15), 
                           DATAIN(14) => data_in(14), DATAIN(13) => data_in(13)
                           , DATAIN(12) => data_in(12), DATAIN(11) => 
                           data_in(11), DATAIN(10) => data_in(10), DATAIN(9) =>
                           data_in(9), DATAIN(8) => data_in(8), DATAIN(7) => 
                           data_in(7), DATAIN(6) => data_in(6), DATAIN(5) => 
                           data_in(5), DATAIN(4) => data_in(4), DATAIN(3) => 
                           data_in(3), DATAIN(2) => data_in(2), DATAIN(1) => 
                           data_in(1), DATAIN(0) => data_in(0), OUT1(63) => 
                           out_1(63), OUT1(62) => out_1(62), OUT1(61) => 
                           out_1(61), OUT1(60) => out_1(60), OUT1(59) => 
                           out_1(59), OUT1(58) => out_1(58), OUT1(57) => 
                           out_1(57), OUT1(56) => out_1(56), OUT1(55) => 
                           out_1(55), OUT1(54) => out_1(54), OUT1(53) => 
                           out_1(53), OUT1(52) => out_1(52), OUT1(51) => 
                           out_1(51), OUT1(50) => out_1(50), OUT1(49) => 
                           out_1(49), OUT1(48) => out_1(48), OUT1(47) => 
                           out_1(47), OUT1(46) => out_1(46), OUT1(45) => 
                           out_1(45), OUT1(44) => out_1(44), OUT1(43) => 
                           out_1(43), OUT1(42) => out_1(42), OUT1(41) => 
                           out_1(41), OUT1(40) => out_1(40), OUT1(39) => 
                           out_1(39), OUT1(38) => out_1(38), OUT1(37) => 
                           out_1(37), OUT1(36) => out_1(36), OUT1(35) => 
                           out_1(35), OUT1(34) => out_1(34), OUT1(33) => 
                           out_1(33), OUT1(32) => out_1(32), OUT1(31) => 
                           out_1(31), OUT1(30) => out_1(30), OUT1(29) => 
                           out_1(29), OUT1(28) => out_1(28), OUT1(27) => 
                           out_1(27), OUT1(26) => out_1(26), OUT1(25) => 
                           out_1(25), OUT1(24) => out_1(24), OUT1(23) => 
                           out_1(23), OUT1(22) => out_1(22), OUT1(21) => 
                           out_1(21), OUT1(20) => out_1(20), OUT1(19) => 
                           out_1(19), OUT1(18) => out_1(18), OUT1(17) => 
                           out_1(17), OUT1(16) => out_1(16), OUT1(15) => 
                           out_1(15), OUT1(14) => out_1(14), OUT1(13) => 
                           out_1(13), OUT1(12) => out_1(12), OUT1(11) => 
                           out_1(11), OUT1(10) => out_1(10), OUT1(9) => 
                           out_1(9), OUT1(8) => out_1(8), OUT1(7) => out_1(7), 
                           OUT1(6) => out_1(6), OUT1(5) => out_1(5), OUT1(4) =>
                           out_1(4), OUT1(3) => out_1(3), OUT1(2) => out_1(2), 
                           OUT1(1) => out_1(1), OUT1(0) => out_1(0), OUT2(63) 
                           => out_2(63), OUT2(62) => out_2(62), OUT2(61) => 
                           out_2(61), OUT2(60) => out_2(60), OUT2(59) => 
                           out_2(59), OUT2(58) => out_2(58), OUT2(57) => 
                           out_2(57), OUT2(56) => out_2(56), OUT2(55) => 
                           out_2(55), OUT2(54) => out_2(54), OUT2(53) => 
                           out_2(53), OUT2(52) => out_2(52), OUT2(51) => 
                           out_2(51), OUT2(50) => out_2(50), OUT2(49) => 
                           out_2(49), OUT2(48) => out_2(48), OUT2(47) => 
                           out_2(47), OUT2(46) => out_2(46), OUT2(45) => 
                           out_2(45), OUT2(44) => out_2(44), OUT2(43) => 
                           out_2(43), OUT2(42) => out_2(42), OUT2(41) => 
                           out_2(41), OUT2(40) => out_2(40), OUT2(39) => 
                           out_2(39), OUT2(38) => out_2(38), OUT2(37) => 
                           out_2(37), OUT2(36) => out_2(36), OUT2(35) => 
                           out_2(35), OUT2(34) => out_2(34), OUT2(33) => 
                           out_2(33), OUT2(32) => out_2(32), OUT2(31) => 
                           out_2(31), OUT2(30) => out_2(30), OUT2(29) => 
                           out_2(29), OUT2(28) => out_2(28), OUT2(27) => 
                           out_2(27), OUT2(26) => out_2(26), OUT2(25) => 
                           out_2(25), OUT2(24) => out_2(24), OUT2(23) => 
                           out_2(23), OUT2(22) => out_2(22), OUT2(21) => 
                           out_2(21), OUT2(20) => out_2(20), OUT2(19) => 
                           out_2(19), OUT2(18) => out_2(18), OUT2(17) => 
                           out_2(17), OUT2(16) => out_2(16), OUT2(15) => 
                           out_2(15), OUT2(14) => out_2(14), OUT2(13) => 
                           out_2(13), OUT2(12) => out_2(12), OUT2(11) => 
                           out_2(11), OUT2(10) => out_2(10), OUT2(9) => 
                           out_2(9), OUT2(8) => out_2(8), OUT2(7) => out_2(7), 
                           OUT2(6) => out_2(6), OUT2(5) => out_2(5), OUT2(4) =>
                           out_2(4), OUT2(3) => out_2(3), OUT2(2) => out_2(2), 
                           OUT2(1) => out_2(1), OUT2(0) => out_2(0));
   r341 : Logix_control_rf_DW01_incdec_0_DW01_incdec_1 port map( A(31) => 
                           cansave_31_port, A(30) => cansave_30_port, A(29) => 
                           cansave_29_port, A(28) => cansave_28_port, A(27) => 
                           cansave_27_port, A(26) => cansave_26_port, A(25) => 
                           cansave_25_port, A(24) => cansave_24_port, A(23) => 
                           cansave_23_port, A(22) => cansave_22_port, A(21) => 
                           cansave_21_port, A(20) => cansave_20_port, A(19) => 
                           cansave_19_port, A(18) => cansave_18_port, A(17) => 
                           cansave_17_port, A(16) => cansave_16_port, A(15) => 
                           cansave_15_port, A(14) => cansave_14_port, A(13) => 
                           cansave_13_port, A(12) => cansave_12_port, A(11) => 
                           cansave_11_port, A(10) => cansave_10_port, A(9) => 
                           cansave_9_port, A(8) => cansave_8_port, A(7) => 
                           cansave_7_port, A(6) => cansave_6_port, A(5) => 
                           cansave_5_port, A(4) => cansave_4_port, A(3) => 
                           cansave_3_port, A(2) => cansave_2_port, A(1) => 
                           cansave_1_port, A(0) => cansave_0_port, INC_DEC => 
                           n867, SUM(31) => N277, SUM(30) => N276, SUM(29) => 
                           N275, SUM(28) => N274, SUM(27) => N273, SUM(26) => 
                           N272, SUM(25) => N271, SUM(24) => N270, SUM(23) => 
                           N269, SUM(22) => N268, SUM(21) => N267, SUM(20) => 
                           N266, SUM(19) => N265, SUM(18) => N264, SUM(17) => 
                           N263, SUM(16) => N262, SUM(15) => N261, SUM(14) => 
                           N260, SUM(13) => N259, SUM(12) => N258, SUM(11) => 
                           N257, SUM(10) => N256, SUM(9) => N255, SUM(8) => 
                           N254, SUM(7) => N253, SUM(6) => N252, SUM(5) => N251
                           , SUM(4) => N250, SUM(3) => N249, SUM(2) => N248, 
                           SUM(1) => N247, SUM(0) => N246);
   r87 : Logix_control_rf_DW01_incdec_1_DW01_incdec_2 port map( A(31) => 
                           canrestore_31_port, A(30) => canrestore_30_port, 
                           A(29) => canrestore_29_port, A(28) => 
                           canrestore_28_port, A(27) => canrestore_27_port, 
                           A(26) => canrestore_26_port, A(25) => 
                           canrestore_25_port, A(24) => canrestore_24_port, 
                           A(23) => canrestore_23_port, A(22) => 
                           canrestore_22_port, A(21) => canrestore_21_port, 
                           A(20) => canrestore_20_port, A(19) => 
                           canrestore_19_port, A(18) => canrestore_18_port, 
                           A(17) => canrestore_17_port, A(16) => 
                           canrestore_16_port, A(15) => canrestore_15_port, 
                           A(14) => canrestore_14_port, A(13) => 
                           canrestore_13_port, A(12) => canrestore_12_port, 
                           A(11) => canrestore_11_port, A(10) => 
                           canrestore_10_port, A(9) => canrestore_9_port, A(8) 
                           => canrestore_8_port, A(7) => canrestore_7_port, 
                           A(6) => canrestore_6_port, A(5) => canrestore_5_port
                           , A(4) => canrestore_4_port, A(3) => 
                           canrestore_3_port, A(2) => canrestore_2_port, A(1) 
                           => canrestore_1_port, A(0) => canrestore_0_port, 
                           INC_DEC => n866, SUM(31) => N676, SUM(30) => N675, 
                           SUM(29) => N674, SUM(28) => N673, SUM(27) => N672, 
                           SUM(26) => N671, SUM(25) => N670, SUM(24) => N669, 
                           SUM(23) => N668, SUM(22) => N667, SUM(21) => N666, 
                           SUM(20) => N665, SUM(19) => N664, SUM(18) => N663, 
                           SUM(17) => N662, SUM(16) => N661, SUM(15) => N660, 
                           SUM(14) => N659, SUM(13) => N658, SUM(12) => N657, 
                           SUM(11) => N656, SUM(10) => N655, SUM(9) => N654, 
                           SUM(8) => N653, SUM(7) => N652, SUM(6) => N651, 
                           SUM(5) => N650, SUM(4) => N649, SUM(3) => N648, 
                           SUM(2) => N647, SUM(1) => N646, SUM(0) => N645);
   memory_bus_tri_0_inst : TBUF_X1 port map( A => n1260, EN => n1259, Z => 
                           memory_bus(0));
   memory_bus_tri_1_inst : TBUF_X1 port map( A => n1133, EN => n1134, Z => 
                           memory_bus(1));
   memory_bus_tri_2_inst : TBUF_X1 port map( A => n1159, EN => n1160, Z => 
                           memory_bus(2));
   memory_bus_tri_3_inst : TBUF_X1 port map( A => n1157, EN => n1158, Z => 
                           memory_bus(3));
   memory_bus_tri_4_inst : TBUF_X1 port map( A => n1155, EN => n1156, Z => 
                           memory_bus(4));
   memory_bus_tri_5_inst : TBUF_X1 port map( A => n1153, EN => n1154, Z => 
                           memory_bus(5));
   memory_bus_tri_6_inst : TBUF_X1 port map( A => n1151, EN => n1152, Z => 
                           memory_bus(6));
   memory_bus_tri_7_inst : TBUF_X1 port map( A => n1149, EN => n1150, Z => 
                           memory_bus(7));
   memory_bus_tri_8_inst : TBUF_X1 port map( A => n1147, EN => n1148, Z => 
                           memory_bus(8));
   memory_bus_tri_9_inst : TBUF_X1 port map( A => n1145, EN => n1146, Z => 
                           memory_bus(9));
   memory_bus_tri_10_inst : TBUF_X1 port map( A => n1143, EN => n1144, Z => 
                           memory_bus(10));
   memory_bus_tri_11_inst : TBUF_X1 port map( A => n1141, EN => n1142, Z => 
                           memory_bus(11));
   memory_bus_tri_12_inst : TBUF_X1 port map( A => n1139, EN => n1140, Z => 
                           memory_bus(12));
   memory_bus_tri_13_inst : TBUF_X1 port map( A => n1137, EN => n1138, Z => 
                           memory_bus(13));
   memory_bus_tri_14_inst : TBUF_X1 port map( A => n1135, EN => n1136, Z => 
                           memory_bus(14));
   memory_bus_tri_15_inst : TBUF_X1 port map( A => n1162, EN => n1161, Z => 
                           memory_bus(15));
   memory_bus_tri_16_inst : TBUF_X1 port map( A => n1164, EN => n1163, Z => 
                           memory_bus(16));
   memory_bus_tri_17_inst : TBUF_X1 port map( A => n1166, EN => n1165, Z => 
                           memory_bus(17));
   memory_bus_tri_18_inst : TBUF_X1 port map( A => n1168, EN => n1167, Z => 
                           memory_bus(18));
   memory_bus_tri_19_inst : TBUF_X1 port map( A => n1170, EN => n1169, Z => 
                           memory_bus(19));
   memory_bus_tri_20_inst : TBUF_X1 port map( A => n1172, EN => n1171, Z => 
                           memory_bus(20));
   memory_bus_tri_21_inst : TBUF_X1 port map( A => n1174, EN => n1173, Z => 
                           memory_bus(21));
   memory_bus_tri_22_inst : TBUF_X1 port map( A => n1176, EN => n1175, Z => 
                           memory_bus(22));
   memory_bus_tri_23_inst : TBUF_X1 port map( A => n1178, EN => n1177, Z => 
                           memory_bus(23));
   memory_bus_tri_24_inst : TBUF_X1 port map( A => n1180, EN => n1179, Z => 
                           memory_bus(24));
   memory_bus_tri_25_inst : TBUF_X1 port map( A => n1182, EN => n1181, Z => 
                           memory_bus(25));
   memory_bus_tri_26_inst : TBUF_X1 port map( A => n1184, EN => n1183, Z => 
                           memory_bus(26));
   memory_bus_tri_27_inst : TBUF_X1 port map( A => n1186, EN => n1185, Z => 
                           memory_bus(27));
   memory_bus_tri_28_inst : TBUF_X1 port map( A => n1188, EN => n1187, Z => 
                           memory_bus(28));
   memory_bus_tri_29_inst : TBUF_X1 port map( A => n1190, EN => n1189, Z => 
                           memory_bus(29));
   memory_bus_tri_30_inst : TBUF_X1 port map( A => n1192, EN => n1191, Z => 
                           memory_bus(30));
   memory_bus_tri_31_inst : TBUF_X1 port map( A => n1194, EN => n1193, Z => 
                           memory_bus(31));
   memory_bus_tri_32_inst : TBUF_X1 port map( A => n1196, EN => n1195, Z => 
                           memory_bus(32));
   memory_bus_tri_33_inst : TBUF_X1 port map( A => n1198, EN => n1197, Z => 
                           memory_bus(33));
   memory_bus_tri_34_inst : TBUF_X1 port map( A => n1200, EN => n1199, Z => 
                           memory_bus(34));
   memory_bus_tri_35_inst : TBUF_X1 port map( A => n1202, EN => n1201, Z => 
                           memory_bus(35));
   memory_bus_tri_36_inst : TBUF_X1 port map( A => n1204, EN => n1203, Z => 
                           memory_bus(36));
   memory_bus_tri_37_inst : TBUF_X1 port map( A => n1206, EN => n1205, Z => 
                           memory_bus(37));
   memory_bus_tri_38_inst : TBUF_X1 port map( A => n1208, EN => n1207, Z => 
                           memory_bus(38));
   memory_bus_tri_39_inst : TBUF_X1 port map( A => n1210, EN => n1209, Z => 
                           memory_bus(39));
   memory_bus_tri_40_inst : TBUF_X1 port map( A => n1212, EN => n1211, Z => 
                           memory_bus(40));
   memory_bus_tri_41_inst : TBUF_X1 port map( A => n1214, EN => n1213, Z => 
                           memory_bus(41));
   memory_bus_tri_42_inst : TBUF_X1 port map( A => n1216, EN => n1215, Z => 
                           memory_bus(42));
   memory_bus_tri_43_inst : TBUF_X1 port map( A => n1218, EN => n1217, Z => 
                           memory_bus(43));
   memory_bus_tri_44_inst : TBUF_X1 port map( A => n1220, EN => n1219, Z => 
                           memory_bus(44));
   memory_bus_tri_45_inst : TBUF_X1 port map( A => n1222, EN => n1221, Z => 
                           memory_bus(45));
   memory_bus_tri_46_inst : TBUF_X1 port map( A => n1224, EN => n1223, Z => 
                           memory_bus(46));
   memory_bus_tri_47_inst : TBUF_X1 port map( A => n1226, EN => n1225, Z => 
                           memory_bus(47));
   memory_bus_tri_48_inst : TBUF_X1 port map( A => n1228, EN => n1227, Z => 
                           memory_bus(48));
   memory_bus_tri_49_inst : TBUF_X1 port map( A => n1230, EN => n1229, Z => 
                           memory_bus(49));
   memory_bus_tri_50_inst : TBUF_X1 port map( A => n1232, EN => n1231, Z => 
                           memory_bus(50));
   memory_bus_tri_51_inst : TBUF_X1 port map( A => n1234, EN => n1233, Z => 
                           memory_bus(51));
   memory_bus_tri_52_inst : TBUF_X1 port map( A => n1236, EN => n1235, Z => 
                           memory_bus(52));
   memory_bus_tri_53_inst : TBUF_X1 port map( A => n1238, EN => n1237, Z => 
                           memory_bus(53));
   memory_bus_tri_54_inst : TBUF_X1 port map( A => n1240, EN => n1239, Z => 
                           memory_bus(54));
   memory_bus_tri_55_inst : TBUF_X1 port map( A => n1242, EN => n1241, Z => 
                           memory_bus(55));
   memory_bus_tri_56_inst : TBUF_X1 port map( A => n1244, EN => n1243, Z => 
                           memory_bus(56));
   memory_bus_tri_57_inst : TBUF_X1 port map( A => n1246, EN => n1245, Z => 
                           memory_bus(57));
   memory_bus_tri_58_inst : TBUF_X1 port map( A => n1248, EN => n1247, Z => 
                           memory_bus(58));
   memory_bus_tri_59_inst : TBUF_X1 port map( A => n1250, EN => n1249, Z => 
                           memory_bus(59));
   memory_bus_tri_60_inst : TBUF_X1 port map( A => n1252, EN => n1251, Z => 
                           memory_bus(60));
   memory_bus_tri_61_inst : TBUF_X1 port map( A => n1254, EN => n1253, Z => 
                           memory_bus(61));
   memory_bus_tri_62_inst : TBUF_X1 port map( A => n1256, EN => n1255, Z => 
                           memory_bus(62));
   memory_bus_tri_63_inst : TBUF_X1 port map( A => n1258, EN => n1257, Z => 
                           memory_bus(63));
   U555 : NOR2_X2 port map( A1 => n975, A2 => n1044, ZN => n864);
   U556 : NOR2_X2 port map( A1 => n975, A2 => n1044, ZN => n865);
   U557 : NOR2_X2 port map( A1 => n975, A2 => n1044, ZN => n976);
   U558 : NAND2_X4 port map( A1 => n972, A2 => n934, ZN => n870);
   U559 : OR2_X4 port map( A1 => n1042, A2 => rest, ZN => n979);
   U560 : NAND2_X4 port map( A1 => n1045, A2 => n878, ZN => n975);
   U561 : AND2_X4 port map( A1 => n978, A2 => n970, ZN => n977);
   U562 : INV_X4 port map( A => n975, ZN => n978);
   U563 : NAND3_X2 port map( A1 => n873, A2 => n964, A3 => n915, ZN => n928);
   U564 : CLKBUF_X3 port map( A => U3_U6_Z_0, Z => n866);
   U565 : NAND3_X2 port map( A1 => n881, A2 => n914, A3 => n915, ZN => n883);
   U566 : INV_X4 port map( A => n918, ZN => n867);
   U567 : BUF_X8 port map( A => clock, Z => n868);
   U568 : BUF_X1 port map( A => clock, Z => n869);
   U569 : OAI22_X1 port map( A1 => n466, A2 => n870, B1 => n871, B2 => n872, ZN
                           => n795);
   U570 : AOI21_X1 port map( B1 => N246, B2 => n873, A => n874, ZN => n871);
   U571 : NAND2_X1 port map( A1 => n875, A2 => n876, ZN => n794);
   U572 : NAND3_X1 port map( A1 => n877, A2 => n878, A3 => n879, ZN => n876);
   U573 : OAI22_X1 port map( A1 => n465, A2 => n870, B1 => n880, B2 => n872, ZN
                           => n793);
   U574 : AOI21_X1 port map( B1 => N645, B2 => n881, A => n882, ZN => n880);
   U575 : OAI22_X1 port map( A1 => n464, A2 => n870, B1 => n883, B2 => n884, ZN
                           => n792);
   U576 : INV_X1 port map( A => N676, ZN => n884);
   U577 : OAI22_X1 port map( A1 => n463, A2 => n870, B1 => n883, B2 => n885, ZN
                           => n791);
   U578 : INV_X1 port map( A => N675, ZN => n885);
   U579 : OAI22_X1 port map( A1 => n462, A2 => n870, B1 => n883, B2 => n886, ZN
                           => n790);
   U580 : INV_X1 port map( A => N674, ZN => n886);
   U581 : OAI22_X1 port map( A1 => n461, A2 => n870, B1 => n883, B2 => n887, ZN
                           => n789);
   U582 : INV_X1 port map( A => N673, ZN => n887);
   U583 : OAI22_X1 port map( A1 => n460, A2 => n870, B1 => n883, B2 => n888, ZN
                           => n788);
   U584 : INV_X1 port map( A => N672, ZN => n888);
   U585 : OAI22_X1 port map( A1 => n459, A2 => n870, B1 => n883, B2 => n889, ZN
                           => n787);
   U586 : INV_X1 port map( A => N671, ZN => n889);
   U587 : OAI22_X1 port map( A1 => n458, A2 => n870, B1 => n883, B2 => n890, ZN
                           => n786);
   U588 : INV_X1 port map( A => N670, ZN => n890);
   U589 : OAI22_X1 port map( A1 => n457, A2 => n870, B1 => n883, B2 => n891, ZN
                           => n785);
   U590 : INV_X1 port map( A => N669, ZN => n891);
   U591 : OAI22_X1 port map( A1 => n456, A2 => n870, B1 => n883, B2 => n892, ZN
                           => n784);
   U592 : INV_X1 port map( A => N668, ZN => n892);
   U593 : OAI22_X1 port map( A1 => n455, A2 => n870, B1 => n883, B2 => n893, ZN
                           => n783);
   U594 : INV_X1 port map( A => N667, ZN => n893);
   U595 : OAI22_X1 port map( A1 => n454, A2 => n870, B1 => n883, B2 => n894, ZN
                           => n782);
   U596 : INV_X1 port map( A => N666, ZN => n894);
   U597 : OAI22_X1 port map( A1 => n453, A2 => n870, B1 => n883, B2 => n895, ZN
                           => n781);
   U598 : INV_X1 port map( A => N665, ZN => n895);
   U599 : OAI22_X1 port map( A1 => n452, A2 => n870, B1 => n883, B2 => n896, ZN
                           => n780);
   U600 : INV_X1 port map( A => N664, ZN => n896);
   U601 : OAI22_X1 port map( A1 => n451, A2 => n870, B1 => n883, B2 => n897, ZN
                           => n779);
   U602 : INV_X1 port map( A => N663, ZN => n897);
   U603 : OAI22_X1 port map( A1 => n450, A2 => n870, B1 => n883, B2 => n898, ZN
                           => n778);
   U604 : INV_X1 port map( A => N662, ZN => n898);
   U605 : OAI22_X1 port map( A1 => n449, A2 => n870, B1 => n883, B2 => n899, ZN
                           => n777);
   U606 : INV_X1 port map( A => N661, ZN => n899);
   U607 : OAI22_X1 port map( A1 => n448, A2 => n870, B1 => n883, B2 => n900, ZN
                           => n776);
   U608 : INV_X1 port map( A => N660, ZN => n900);
   U609 : OAI22_X1 port map( A1 => n447, A2 => n870, B1 => n883, B2 => n901, ZN
                           => n775);
   U610 : INV_X1 port map( A => N659, ZN => n901);
   U611 : OAI22_X1 port map( A1 => n446, A2 => n870, B1 => n883, B2 => n902, ZN
                           => n774);
   U612 : INV_X1 port map( A => N658, ZN => n902);
   U613 : OAI22_X1 port map( A1 => n445, A2 => n870, B1 => n883, B2 => n903, ZN
                           => n773);
   U614 : INV_X1 port map( A => N657, ZN => n903);
   U615 : OAI22_X1 port map( A1 => n444, A2 => n870, B1 => n883, B2 => n904, ZN
                           => n772);
   U616 : INV_X1 port map( A => N656, ZN => n904);
   U617 : OAI22_X1 port map( A1 => n443, A2 => n870, B1 => n883, B2 => n905, ZN
                           => n771);
   U618 : INV_X1 port map( A => N655, ZN => n905);
   U619 : OAI22_X1 port map( A1 => n442, A2 => n870, B1 => n883, B2 => n906, ZN
                           => n770);
   U620 : INV_X1 port map( A => N654, ZN => n906);
   U621 : OAI22_X1 port map( A1 => n441, A2 => n870, B1 => n883, B2 => n907, ZN
                           => n769);
   U622 : INV_X1 port map( A => N653, ZN => n907);
   U623 : OAI22_X1 port map( A1 => n440, A2 => n870, B1 => n883, B2 => n908, ZN
                           => n768);
   U624 : INV_X1 port map( A => N652, ZN => n908);
   U625 : OAI22_X1 port map( A1 => n439, A2 => n870, B1 => n883, B2 => n909, ZN
                           => n767);
   U626 : INV_X1 port map( A => N651, ZN => n909);
   U627 : OAI22_X1 port map( A1 => n438, A2 => n870, B1 => n883, B2 => n910, ZN
                           => n766);
   U628 : INV_X1 port map( A => N650, ZN => n910);
   U629 : OAI22_X1 port map( A1 => n437, A2 => n870, B1 => n883, B2 => n911, ZN
                           => n765);
   U630 : INV_X1 port map( A => N649, ZN => n911);
   U631 : OAI22_X1 port map( A1 => n436, A2 => n870, B1 => n883, B2 => n912, ZN
                           => n764);
   U632 : INV_X1 port map( A => N648, ZN => n912);
   U633 : OAI22_X1 port map( A1 => n435, A2 => n870, B1 => n883, B2 => n913, ZN
                           => n763);
   U634 : INV_X1 port map( A => N647, ZN => n913);
   U635 : INV_X1 port map( A => n882, ZN => n914);
   U636 : OAI22_X1 port map( A1 => n434, A2 => n870, B1 => n916, B2 => n872, ZN
                           => n762);
   U637 : AOI21_X1 port map( B1 => N646, B2 => n881, A => n882, ZN => n916);
   U638 : NOR2_X1 port map( A1 => n917, A2 => n918, ZN => n882);
   U639 : NAND2_X1 port map( A1 => n918, A2 => n917, ZN => n881);
   U640 : NAND2_X1 port map( A1 => n464, A2 => n919, ZN => n917);
   U641 : OAI221_X1 port map( B1 => n465, B2 => n434, C1 => r339_LEQ, C2 => 
                           n920, A => n921, ZN => n919);
   U642 : MUX2_X1 port map( A => N1274, B => n922, S => n923, Z => n761);
   U643 : INV_X1 port map( A => n924, ZN => n922);
   U644 : AOI22_X1 port map( A1 => n925, A2 => n433, B1 => n878, B2 => n926, ZN
                           => n924);
   U645 : OAI22_X1 port map( A1 => n432, A2 => n870, B1 => n927, B2 => n872, ZN
                           => n760);
   U646 : AOI21_X1 port map( B1 => N247, B2 => n873, A => n874, ZN => n927);
   U647 : OAI22_X1 port map( A1 => n431, A2 => n870, B1 => n928, B2 => n929, ZN
                           => n759);
   U648 : INV_X1 port map( A => N277, ZN => n929);
   U649 : MUX2_X1 port map( A => n930, B => cansave_2_port, S => n931, Z => 
                           n758);
   U650 : OAI21_X1 port map( B1 => n932, B2 => n933, A => n934, ZN => n930);
   U651 : XOR2_X1 port map( A => n918, B => n935, Z => n933);
   U652 : INV_X1 port map( A => r339_LEQ, ZN => n918);
   U653 : INV_X1 port map( A => N248, ZN => n932);
   U654 : OAI22_X1 port map( A1 => n429, A2 => n870, B1 => n928, B2 => n936, ZN
                           => n757);
   U655 : INV_X1 port map( A => N276, ZN => n936);
   U656 : OAI22_X1 port map( A1 => n428, A2 => n870, B1 => n928, B2 => n937, ZN
                           => n756);
   U657 : INV_X1 port map( A => N275, ZN => n937);
   U658 : OAI22_X1 port map( A1 => n427, A2 => n870, B1 => n928, B2 => n938, ZN
                           => n755);
   U659 : INV_X1 port map( A => N274, ZN => n938);
   U660 : OAI22_X1 port map( A1 => n426, A2 => n870, B1 => n928, B2 => n939, ZN
                           => n754);
   U661 : INV_X1 port map( A => N273, ZN => n939);
   U662 : OAI22_X1 port map( A1 => n425, A2 => n870, B1 => n928, B2 => n940, ZN
                           => n753);
   U663 : INV_X1 port map( A => N272, ZN => n940);
   U664 : OAI22_X1 port map( A1 => n424, A2 => n870, B1 => n928, B2 => n941, ZN
                           => n752);
   U665 : INV_X1 port map( A => N271, ZN => n941);
   U666 : OAI22_X1 port map( A1 => n423, A2 => n870, B1 => n928, B2 => n942, ZN
                           => n751);
   U667 : INV_X1 port map( A => N270, ZN => n942);
   U668 : OAI22_X1 port map( A1 => n422, A2 => n870, B1 => n928, B2 => n943, ZN
                           => n750);
   U669 : INV_X1 port map( A => N269, ZN => n943);
   U670 : OAI22_X1 port map( A1 => n421, A2 => n870, B1 => n928, B2 => n944, ZN
                           => n749);
   U671 : INV_X1 port map( A => N268, ZN => n944);
   U672 : OAI22_X1 port map( A1 => n420, A2 => n870, B1 => n928, B2 => n945, ZN
                           => n748);
   U673 : INV_X1 port map( A => N267, ZN => n945);
   U674 : OAI22_X1 port map( A1 => n419, A2 => n870, B1 => n928, B2 => n946, ZN
                           => n747);
   U675 : INV_X1 port map( A => N266, ZN => n946);
   U676 : OAI22_X1 port map( A1 => n418, A2 => n870, B1 => n928, B2 => n947, ZN
                           => n746);
   U677 : INV_X1 port map( A => N265, ZN => n947);
   U678 : OAI22_X1 port map( A1 => n417, A2 => n870, B1 => n928, B2 => n948, ZN
                           => n745);
   U679 : INV_X1 port map( A => N264, ZN => n948);
   U680 : OAI22_X1 port map( A1 => n416, A2 => n870, B1 => n928, B2 => n949, ZN
                           => n744);
   U681 : INV_X1 port map( A => N263, ZN => n949);
   U682 : OAI22_X1 port map( A1 => n415, A2 => n870, B1 => n928, B2 => n950, ZN
                           => n743);
   U683 : INV_X1 port map( A => N262, ZN => n950);
   U684 : OAI22_X1 port map( A1 => n414, A2 => n870, B1 => n928, B2 => n951, ZN
                           => n742);
   U685 : INV_X1 port map( A => N261, ZN => n951);
   U686 : OAI22_X1 port map( A1 => n413, A2 => n870, B1 => n928, B2 => n952, ZN
                           => n741);
   U687 : INV_X1 port map( A => N260, ZN => n952);
   U688 : OAI22_X1 port map( A1 => n412, A2 => n870, B1 => n928, B2 => n953, ZN
                           => n740);
   U689 : INV_X1 port map( A => N259, ZN => n953);
   U690 : OAI22_X1 port map( A1 => n411, A2 => n870, B1 => n928, B2 => n954, ZN
                           => n739);
   U691 : INV_X1 port map( A => N258, ZN => n954);
   U692 : OAI22_X1 port map( A1 => n410, A2 => n870, B1 => n928, B2 => n955, ZN
                           => n738);
   U693 : INV_X1 port map( A => N257, ZN => n955);
   U694 : OAI22_X1 port map( A1 => n409, A2 => n870, B1 => n928, B2 => n956, ZN
                           => n737);
   U695 : INV_X1 port map( A => N256, ZN => n956);
   U696 : OAI22_X1 port map( A1 => n408, A2 => n870, B1 => n928, B2 => n957, ZN
                           => n736);
   U697 : INV_X1 port map( A => N255, ZN => n957);
   U698 : OAI22_X1 port map( A1 => n407, A2 => n870, B1 => n928, B2 => n958, ZN
                           => n735);
   U699 : INV_X1 port map( A => N254, ZN => n958);
   U700 : OAI22_X1 port map( A1 => n406, A2 => n870, B1 => n928, B2 => n959, ZN
                           => n734);
   U701 : INV_X1 port map( A => N253, ZN => n959);
   U702 : OAI22_X1 port map( A1 => n405, A2 => n870, B1 => n928, B2 => n960, ZN
                           => n733);
   U703 : INV_X1 port map( A => N252, ZN => n960);
   U704 : OAI22_X1 port map( A1 => n404, A2 => n870, B1 => n928, B2 => n961, ZN
                           => n732);
   U705 : INV_X1 port map( A => N251, ZN => n961);
   U706 : OAI22_X1 port map( A1 => n403, A2 => n870, B1 => n928, B2 => n962, ZN
                           => n731);
   U707 : INV_X1 port map( A => N250, ZN => n962);
   U708 : OAI22_X1 port map( A1 => n402, A2 => n870, B1 => n928, B2 => n963, ZN
                           => n730);
   U709 : INV_X1 port map( A => N249, ZN => n963);
   U710 : INV_X1 port map( A => n872, ZN => n915);
   U711 : NAND2_X1 port map( A1 => n925, A2 => n870, ZN => n872);
   U712 : INV_X1 port map( A => n874, ZN => n964);
   U713 : NOR2_X1 port map( A1 => n935, A2 => r339_LEQ, ZN => n874);
   U714 : NAND2_X1 port map( A1 => r339_LEQ, A2 => n935, ZN => n873);
   U715 : NAND2_X1 port map( A1 => n431, A2 => n965, ZN => n935);
   U716 : OAI211_X1 port map( C1 => n466, C2 => n432, A => n866, B => n966, ZN 
                           => n965);
   U717 : AOI21_X1 port map( B1 => n931, B2 => n1130, A => n967, ZN => n729);
   U718 : AOI22_X1 port map( A1 => n968, A2 => n969, B1 => n970, B2 => n878, ZN
                           => n967);
   U719 : NOR2_X1 port map( A1 => call, A2 => n971, ZN => n968);
   U720 : INV_X1 port map( A => n870, ZN => n931);
   U721 : OAI21_X1 port map( B1 => ret, B2 => call, A => n973, ZN => n972);
   U722 : INV_X1 port map( A => n974, ZN => n728);
   U723 : AOI221_X1 port map( B1 => n1133, B2 => n975, C1 => data_in(1), C2 => 
                           n976, A => n977, ZN => n974);
   U724 : OAI21_X1 port map( B1 => n978, B2 => n829, A => n979, ZN => n727);
   U725 : INV_X1 port map( A => n980, ZN => n726);
   U726 : AOI221_X1 port map( B1 => n1135, B2 => n975, C1 => data_in(14), C2 =>
                           n865, A => n977, ZN => n980);
   U727 : OAI21_X1 port map( B1 => n978, B2 => n830, A => n979, ZN => n725);
   U728 : INV_X1 port map( A => n981, ZN => n724);
   U729 : AOI221_X1 port map( B1 => n1137, B2 => n975, C1 => data_in(13), C2 =>
                           n864, A => n977, ZN => n981);
   U730 : OAI21_X1 port map( B1 => n978, B2 => n831, A => n979, ZN => n723);
   U731 : INV_X1 port map( A => n982, ZN => n722);
   U732 : AOI221_X1 port map( B1 => n1139, B2 => n975, C1 => data_in(12), C2 =>
                           n976, A => n977, ZN => n982);
   U733 : OAI21_X1 port map( B1 => n978, B2 => n832, A => n979, ZN => n721);
   U734 : INV_X1 port map( A => n983, ZN => n720);
   U735 : AOI221_X1 port map( B1 => n1141, B2 => n975, C1 => data_in(11), C2 =>
                           n865, A => n977, ZN => n983);
   U736 : OAI21_X1 port map( B1 => n978, B2 => n833, A => n979, ZN => n719);
   U737 : INV_X1 port map( A => n984, ZN => n718);
   U738 : AOI221_X1 port map( B1 => n1143, B2 => n975, C1 => data_in(10), C2 =>
                           n864, A => n977, ZN => n984);
   U739 : OAI21_X1 port map( B1 => n978, B2 => n834, A => n979, ZN => n717);
   U740 : INV_X1 port map( A => n985, ZN => n716);
   U741 : AOI221_X1 port map( B1 => n1145, B2 => n975, C1 => data_in(9), C2 => 
                           n976, A => n977, ZN => n985);
   U742 : OAI21_X1 port map( B1 => n978, B2 => n835, A => n979, ZN => n715);
   U743 : INV_X1 port map( A => n986, ZN => n714);
   U744 : AOI221_X1 port map( B1 => n1147, B2 => n975, C1 => data_in(8), C2 => 
                           n865, A => n977, ZN => n986);
   U745 : OAI21_X1 port map( B1 => n978, B2 => n836, A => n979, ZN => n713);
   U746 : INV_X1 port map( A => n987, ZN => n712);
   U747 : AOI221_X1 port map( B1 => n1149, B2 => n975, C1 => data_in(7), C2 => 
                           n864, A => n977, ZN => n987);
   U748 : OAI21_X1 port map( B1 => n978, B2 => n837, A => n979, ZN => n711);
   U749 : INV_X1 port map( A => n988, ZN => n710);
   U750 : AOI221_X1 port map( B1 => n1151, B2 => n975, C1 => data_in(6), C2 => 
                           n976, A => n977, ZN => n988);
   U751 : OAI21_X1 port map( B1 => n978, B2 => n838, A => n979, ZN => n709);
   U752 : INV_X1 port map( A => n989, ZN => n708);
   U753 : AOI221_X1 port map( B1 => n1153, B2 => n975, C1 => data_in(5), C2 => 
                           n865, A => n977, ZN => n989);
   U754 : OAI21_X1 port map( B1 => n978, B2 => n839, A => n979, ZN => n707);
   U755 : INV_X1 port map( A => n990, ZN => n706);
   U756 : AOI221_X1 port map( B1 => n1155, B2 => n975, C1 => data_in(4), C2 => 
                           n864, A => n977, ZN => n990);
   U757 : OAI21_X1 port map( B1 => n978, B2 => n840, A => n979, ZN => n705);
   U758 : INV_X1 port map( A => n991, ZN => n704);
   U759 : AOI221_X1 port map( B1 => n1157, B2 => n975, C1 => data_in(3), C2 => 
                           n976, A => n977, ZN => n991);
   U760 : OAI21_X1 port map( B1 => n978, B2 => n841, A => n979, ZN => n703);
   U761 : INV_X1 port map( A => n992, ZN => n702);
   U762 : AOI221_X1 port map( B1 => n1159, B2 => n975, C1 => data_in(2), C2 => 
                           n865, A => n977, ZN => n992);
   U763 : OAI21_X1 port map( B1 => n978, B2 => n842, A => n979, ZN => n701);
   U764 : OAI21_X1 port map( B1 => n978, B2 => n843, A => n979, ZN => n700);
   U765 : INV_X1 port map( A => n993, ZN => n699);
   U766 : AOI221_X1 port map( B1 => n1162, B2 => n975, C1 => data_in(15), C2 =>
                           n864, A => n977, ZN => n993);
   U767 : OAI21_X1 port map( B1 => n978, B2 => n844, A => n979, ZN => n698);
   U768 : INV_X1 port map( A => n994, ZN => n697);
   U769 : AOI221_X1 port map( B1 => n1164, B2 => n975, C1 => data_in(16), C2 =>
                           n976, A => n977, ZN => n994);
   U770 : OAI21_X1 port map( B1 => n978, B2 => n845, A => n979, ZN => n696);
   U771 : INV_X1 port map( A => n995, ZN => n695);
   U772 : AOI221_X1 port map( B1 => n1166, B2 => n975, C1 => data_in(17), C2 =>
                           n865, A => n977, ZN => n995);
   U773 : OAI21_X1 port map( B1 => n978, B2 => n846, A => n979, ZN => n694);
   U774 : INV_X1 port map( A => n996, ZN => n693);
   U775 : AOI221_X1 port map( B1 => n1168, B2 => n975, C1 => data_in(18), C2 =>
                           n864, A => n977, ZN => n996);
   U776 : OAI21_X1 port map( B1 => n978, B2 => n847, A => n979, ZN => n692);
   U777 : INV_X1 port map( A => n997, ZN => n691);
   U778 : AOI221_X1 port map( B1 => n1170, B2 => n975, C1 => data_in(19), C2 =>
                           n976, A => n977, ZN => n997);
   U779 : OAI21_X1 port map( B1 => n978, B2 => n848, A => n979, ZN => n690);
   U780 : INV_X1 port map( A => n998, ZN => n689);
   U781 : AOI221_X1 port map( B1 => n1172, B2 => n975, C1 => data_in(20), C2 =>
                           n865, A => n977, ZN => n998);
   U782 : OAI21_X1 port map( B1 => n978, B2 => n849, A => n979, ZN => n688);
   U783 : INV_X1 port map( A => n999, ZN => n687);
   U784 : AOI221_X1 port map( B1 => n1174, B2 => n975, C1 => data_in(21), C2 =>
                           n864, A => n977, ZN => n999);
   U785 : OAI21_X1 port map( B1 => n978, B2 => n850, A => n979, ZN => n686);
   U786 : INV_X1 port map( A => n1000, ZN => n685);
   U787 : AOI221_X1 port map( B1 => n1176, B2 => n975, C1 => data_in(22), C2 =>
                           n976, A => n977, ZN => n1000);
   U788 : OAI21_X1 port map( B1 => n978, B2 => n851, A => n979, ZN => n684);
   U789 : INV_X1 port map( A => n1001, ZN => n683);
   U790 : AOI221_X1 port map( B1 => n1178, B2 => n975, C1 => data_in(23), C2 =>
                           n865, A => n977, ZN => n1001);
   U791 : OAI21_X1 port map( B1 => n978, B2 => n852, A => n979, ZN => n682);
   U792 : INV_X1 port map( A => n1002, ZN => n681);
   U793 : AOI221_X1 port map( B1 => n1180, B2 => n975, C1 => data_in(24), C2 =>
                           n864, A => n977, ZN => n1002);
   U794 : OAI21_X1 port map( B1 => n978, B2 => n853, A => n979, ZN => n680);
   U795 : INV_X1 port map( A => n1003, ZN => n679);
   U796 : AOI221_X1 port map( B1 => n1182, B2 => n975, C1 => data_in(25), C2 =>
                           n976, A => n977, ZN => n1003);
   U797 : OAI21_X1 port map( B1 => n978, B2 => n854, A => n979, ZN => n678);
   U798 : INV_X1 port map( A => n1004, ZN => n677);
   U799 : AOI221_X1 port map( B1 => n1184, B2 => n975, C1 => data_in(26), C2 =>
                           n865, A => n977, ZN => n1004);
   U800 : OAI21_X1 port map( B1 => n978, B2 => n855, A => n979, ZN => n676_port
                           );
   U801 : INV_X1 port map( A => n1005, ZN => n675_port);
   U802 : AOI221_X1 port map( B1 => n1186, B2 => n975, C1 => data_in(27), C2 =>
                           n864, A => n977, ZN => n1005);
   U803 : OAI21_X1 port map( B1 => n978, B2 => n856, A => n979, ZN => n674_port
                           );
   U804 : INV_X1 port map( A => n1006_port, ZN => n673_port);
   U805 : AOI221_X1 port map( B1 => n1188, B2 => n975, C1 => data_in(28), C2 =>
                           n976, A => n977, ZN => n1006_port);
   U806 : OAI21_X1 port map( B1 => n978, B2 => n857, A => n979, ZN => n672_port
                           );
   U807 : INV_X1 port map( A => n1007, ZN => n671_port);
   U808 : AOI221_X1 port map( B1 => n1190, B2 => n975, C1 => data_in(29), C2 =>
                           n865, A => n977, ZN => n1007);
   U809 : OAI21_X1 port map( B1 => n978, B2 => n858, A => n979, ZN => n670_port
                           );
   U810 : INV_X1 port map( A => n1008, ZN => n669_port);
   U811 : AOI221_X1 port map( B1 => n1192, B2 => n975, C1 => data_in(30), C2 =>
                           n864, A => n977, ZN => n1008);
   U812 : OAI21_X1 port map( B1 => n978, B2 => n859, A => n979, ZN => n668_port
                           );
   U813 : INV_X1 port map( A => n1009, ZN => n667_port);
   U814 : AOI221_X1 port map( B1 => n1194, B2 => n975, C1 => data_in(31), C2 =>
                           n976, A => n977, ZN => n1009);
   U815 : OAI21_X1 port map( B1 => n978, B2 => n860, A => n979, ZN => n666_port
                           );
   U816 : INV_X1 port map( A => n1010, ZN => n665_port);
   U817 : AOI221_X1 port map( B1 => n1196, B2 => n975, C1 => data_in(32), C2 =>
                           n865, A => n977, ZN => n1010);
   U818 : OAI21_X1 port map( B1 => n978, B2 => n861, A => n979, ZN => n664_port
                           );
   U819 : INV_X1 port map( A => n1011, ZN => n663_port);
   U820 : AOI221_X1 port map( B1 => n1198, B2 => n975, C1 => data_in(33), C2 =>
                           n864, A => n977, ZN => n1011);
   U821 : OAI21_X1 port map( B1 => n978, B2 => n862, A => n979, ZN => n662_port
                           );
   U822 : INV_X1 port map( A => n1012, ZN => n661_port);
   U823 : AOI221_X1 port map( B1 => n1200, B2 => n975, C1 => data_in(34), C2 =>
                           n976, A => n977, ZN => n1012);
   U824 : OAI21_X1 port map( B1 => n978, B2 => n863, A => n979, ZN => n660_port
                           );
   U825 : INV_X1 port map( A => n1013, ZN => n659_port);
   U826 : AOI221_X1 port map( B1 => n1202, B2 => n975, C1 => data_in(35), C2 =>
                           n865, A => n977, ZN => n1013);
   U827 : OAI21_X1 port map( B1 => n978, B2 => n800, A => n979, ZN => n658_port
                           );
   U828 : INV_X1 port map( A => n1014, ZN => n657_port);
   U829 : AOI221_X1 port map( B1 => n1204, B2 => n975, C1 => data_in(36), C2 =>
                           n864, A => n977, ZN => n1014);
   U830 : OAI21_X1 port map( B1 => n978, B2 => n801, A => n979, ZN => n656_port
                           );
   U831 : INV_X1 port map( A => n1015, ZN => n655_port);
   U832 : AOI221_X1 port map( B1 => n1206, B2 => n975, C1 => data_in(37), C2 =>
                           n976, A => n977, ZN => n1015);
   U833 : OAI21_X1 port map( B1 => n978, B2 => n802, A => n979, ZN => n654_port
                           );
   U834 : INV_X1 port map( A => n1016, ZN => n653_port);
   U835 : AOI221_X1 port map( B1 => n1208, B2 => n975, C1 => data_in(38), C2 =>
                           n865, A => n977, ZN => n1016);
   U836 : OAI21_X1 port map( B1 => n978, B2 => n803, A => n979, ZN => n652_port
                           );
   U837 : INV_X1 port map( A => n1017, ZN => n651_port);
   U838 : AOI221_X1 port map( B1 => n1210, B2 => n975, C1 => data_in(39), C2 =>
                           n864, A => n977, ZN => n1017);
   U839 : OAI21_X1 port map( B1 => n978, B2 => n804, A => n979, ZN => n650_port
                           );
   U840 : INV_X1 port map( A => n1018, ZN => n649_port);
   U841 : AOI221_X1 port map( B1 => n1212, B2 => n975, C1 => data_in(40), C2 =>
                           n976, A => n977, ZN => n1018);
   U842 : OAI21_X1 port map( B1 => n978, B2 => n805, A => n979, ZN => n648_port
                           );
   U843 : INV_X1 port map( A => n1019, ZN => n647_port);
   U844 : AOI221_X1 port map( B1 => n1214, B2 => n975, C1 => data_in(41), C2 =>
                           n865, A => n977, ZN => n1019);
   U845 : OAI21_X1 port map( B1 => n978, B2 => n806, A => n979, ZN => n646_port
                           );
   U846 : INV_X1 port map( A => n1020, ZN => n645_port);
   U847 : AOI221_X1 port map( B1 => n1216, B2 => n975, C1 => data_in(42), C2 =>
                           n864, A => n977, ZN => n1020);
   U848 : OAI21_X1 port map( B1 => n978, B2 => n807, A => n979, ZN => n644);
   U849 : INV_X1 port map( A => n1021, ZN => n643);
   U850 : AOI221_X1 port map( B1 => n1218, B2 => n975, C1 => data_in(43), C2 =>
                           n976, A => n977, ZN => n1021);
   U851 : OAI21_X1 port map( B1 => n978, B2 => n808, A => n979, ZN => n642);
   U852 : INV_X1 port map( A => n1022, ZN => n641);
   U853 : AOI221_X1 port map( B1 => n1220, B2 => n975, C1 => data_in(44), C2 =>
                           n865, A => n977, ZN => n1022);
   U854 : OAI21_X1 port map( B1 => n978, B2 => n809, A => n979, ZN => n640);
   U855 : INV_X1 port map( A => n1023, ZN => n639);
   U856 : AOI221_X1 port map( B1 => n1222, B2 => n975, C1 => data_in(45), C2 =>
                           n864, A => n977, ZN => n1023);
   U857 : OAI21_X1 port map( B1 => n978, B2 => n810, A => n979, ZN => n638);
   U858 : INV_X1 port map( A => n1024, ZN => n637);
   U859 : AOI221_X1 port map( B1 => n1224, B2 => n975, C1 => data_in(46), C2 =>
                           n976, A => n977, ZN => n1024);
   U860 : OAI21_X1 port map( B1 => n978, B2 => n811, A => n979, ZN => n636);
   U861 : INV_X1 port map( A => n1025, ZN => n635);
   U862 : AOI221_X1 port map( B1 => n1226, B2 => n975, C1 => data_in(47), C2 =>
                           n865, A => n977, ZN => n1025);
   U863 : OAI21_X1 port map( B1 => n978, B2 => n812, A => n979, ZN => n634);
   U864 : INV_X1 port map( A => n1026, ZN => n633);
   U865 : AOI221_X1 port map( B1 => n1228, B2 => n975, C1 => data_in(48), C2 =>
                           n864, A => n977, ZN => n1026);
   U866 : OAI21_X1 port map( B1 => n978, B2 => n813, A => n979, ZN => n632);
   U867 : INV_X1 port map( A => n1027, ZN => n631);
   U868 : AOI221_X1 port map( B1 => n1230, B2 => n975, C1 => data_in(49), C2 =>
                           n976, A => n977, ZN => n1027);
   U869 : OAI21_X1 port map( B1 => n978, B2 => n814, A => n979, ZN => n630);
   U870 : INV_X1 port map( A => n1028, ZN => n629);
   U871 : AOI221_X1 port map( B1 => n1232, B2 => n975, C1 => data_in(50), C2 =>
                           n865, A => n977, ZN => n1028);
   U872 : OAI21_X1 port map( B1 => n978, B2 => n815, A => n979, ZN => n628);
   U873 : INV_X1 port map( A => n1029, ZN => n627);
   U874 : AOI221_X1 port map( B1 => n1234, B2 => n975, C1 => data_in(51), C2 =>
                           n864, A => n977, ZN => n1029);
   U875 : OAI21_X1 port map( B1 => n978, B2 => n816, A => n979, ZN => n626);
   U876 : INV_X1 port map( A => n1030, ZN => n625);
   U877 : AOI221_X1 port map( B1 => n1236, B2 => n975, C1 => data_in(52), C2 =>
                           n976, A => n977, ZN => n1030);
   U878 : OAI21_X1 port map( B1 => n978, B2 => n817, A => n979, ZN => n624);
   U879 : INV_X1 port map( A => n1031, ZN => n623);
   U880 : AOI221_X1 port map( B1 => n1238, B2 => n975, C1 => data_in(53), C2 =>
                           n865, A => n977, ZN => n1031);
   U881 : OAI21_X1 port map( B1 => n978, B2 => n818, A => n979, ZN => n622);
   U882 : INV_X1 port map( A => n1032, ZN => n621);
   U883 : AOI221_X1 port map( B1 => n1240, B2 => n975, C1 => data_in(54), C2 =>
                           n864, A => n977, ZN => n1032);
   U884 : OAI21_X1 port map( B1 => n978, B2 => n819, A => n979, ZN => n620);
   U885 : INV_X1 port map( A => n1033, ZN => n619);
   U886 : AOI221_X1 port map( B1 => n1242, B2 => n975, C1 => data_in(55), C2 =>
                           n976, A => n977, ZN => n1033);
   U887 : OAI21_X1 port map( B1 => n978, B2 => n820, A => n979, ZN => n618);
   U888 : INV_X1 port map( A => n1034, ZN => n617);
   U889 : AOI221_X1 port map( B1 => n1244, B2 => n975, C1 => data_in(56), C2 =>
                           n865, A => n977, ZN => n1034);
   U890 : OAI21_X1 port map( B1 => n978, B2 => n821, A => n979, ZN => n616);
   U891 : INV_X1 port map( A => n1035, ZN => n615);
   U892 : AOI221_X1 port map( B1 => n1246, B2 => n975, C1 => data_in(57), C2 =>
                           n864, A => n977, ZN => n1035);
   U893 : OAI21_X1 port map( B1 => n978, B2 => n822, A => n979, ZN => n614);
   U894 : INV_X1 port map( A => n1036, ZN => n613);
   U895 : AOI221_X1 port map( B1 => n1248, B2 => n975, C1 => data_in(58), C2 =>
                           n976, A => n977, ZN => n1036);
   U896 : OAI21_X1 port map( B1 => n978, B2 => n823, A => n979, ZN => n612);
   U897 : INV_X1 port map( A => n1037, ZN => n611);
   U898 : AOI221_X1 port map( B1 => n1250, B2 => n975, C1 => data_in(59), C2 =>
                           n865, A => n977, ZN => n1037);
   U899 : OAI21_X1 port map( B1 => n978, B2 => n824, A => n979, ZN => n610);
   U900 : INV_X1 port map( A => n1038, ZN => n609);
   U901 : AOI221_X1 port map( B1 => n1252, B2 => n975, C1 => data_in(60), C2 =>
                           n864, A => n977, ZN => n1038);
   U902 : OAI21_X1 port map( B1 => n978, B2 => n825, A => n979, ZN => n608);
   U903 : INV_X1 port map( A => n1039, ZN => n607);
   U904 : AOI221_X1 port map( B1 => n1254, B2 => n975, C1 => data_in(61), C2 =>
                           n976, A => n977, ZN => n1039);
   U905 : OAI21_X1 port map( B1 => n978, B2 => n826, A => n979, ZN => n606);
   U906 : INV_X1 port map( A => n1040, ZN => n605);
   U907 : AOI221_X1 port map( B1 => n1256, B2 => n975, C1 => data_in(62), C2 =>
                           n865, A => n977, ZN => n1040);
   U908 : OAI21_X1 port map( B1 => n978, B2 => n827, A => n979, ZN => n604);
   U909 : INV_X1 port map( A => n1041, ZN => n603);
   U910 : AOI221_X1 port map( B1 => n1258, B2 => n975, C1 => data_in(63), C2 =>
                           n864, A => n977, ZN => n1041);
   U911 : OAI21_X1 port map( B1 => n978, B2 => n828, A => n979, ZN => n602);
   U912 : INV_X1 port map( A => n1043, ZN => n601);
   U913 : AOI221_X1 port map( B1 => n1260, B2 => n975, C1 => data_in(0), C2 => 
                           n976, A => n977, ZN => n1043);
   U914 : NOR3_X1 port map( A1 => memory_response, A2 => n1130, A3 => n926, ZN 
                           => n970);
   U915 : OAI21_X1 port map( B1 => n1130, B2 => n926, A => n1044, ZN => n1045);
   U916 : NAND2_X1 port map( A1 => n1046, A2 => n934, ZN => n600);
   U917 : XOR2_X1 port map( A => cwp_o_1_port, B => n1047, Z => n1046);
   U918 : NAND2_X1 port map( A1 => n1048, A2 => n923, ZN => n1047);
   U919 : OAI21_X1 port map( B1 => n1049, B2 => n1050, A => n934, ZN => n923);
   U920 : INV_X1 port map( A => n973, ZN => n1050);
   U921 : NOR2_X1 port map( A1 => r339_LEQ, A2 => n1051, ZN => n1049);
   U922 : NOR2_X1 port map( A1 => n1052, A2 => n1053, ZN => r339_LEQ);
   U923 : XOR2_X1 port map( A => N1274, B => n1051, Z => n1048);
   U924 : AND3_X1 port map( A1 => n1054, A2 => n1052, A3 => ret, ZN => n1051);
   U925 : NAND2_X1 port map( A1 => n875, A2 => n1055, ZN => n599);
   U926 : NAND3_X1 port map( A1 => n1042, A2 => n934, A3 => spill_port, ZN => 
                           n1055);
   U927 : NAND2_X1 port map( A1 => memory_response, A2 => n879, ZN => n1042);
   U928 : NAND3_X1 port map( A1 => n925, A2 => call, A3 => n1053, ZN => n875);
   U929 : NAND2_X1 port map( A1 => n1056, A2 => n1057, ZN => n598);
   U930 : NAND4_X1 port map( A1 => n969, A2 => ret, A3 => n925, A4 => n1052, ZN
                           => n1057);
   U931 : INV_X1 port map( A => n971, ZN => n925);
   U932 : NAND2_X1 port map( A1 => n973, A2 => n878, ZN => n971);
   U933 : INV_X1 port map( A => rest, ZN => n878);
   U934 : NOR2_X1 port map( A1 => n799, A2 => n926, ZN => n973);
   U935 : INV_X1 port map( A => n1054, ZN => n969);
   U936 : NAND3_X1 port map( A1 => n464, A2 => n921, A3 => n920, ZN => n1054);
   U937 : AND2_X1 port map( A1 => n465, A2 => n434, ZN => n920);
   U938 : AND4_X1 port map( A1 => n1058, A2 => n1059, A3 => n1060, A4 => n1061,
                           ZN => n921);
   U939 : NOR2_X1 port map( A1 => n1062, A2 => n1063, ZN => n1061);
   U940 : NAND4_X1 port map( A1 => n442, A2 => n441, A3 => n440, A4 => n439, ZN
                           => n1063);
   U941 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => n1062);
   U942 : AND4_X1 port map( A1 => n1064, A2 => n449, A3 => n447, A4 => n448, ZN
                           => n1060);
   U943 : AND4_X1 port map( A1 => n446, A2 => n445, A3 => n444, A4 => n443, ZN 
                           => n1064);
   U944 : AND4_X1 port map( A1 => n1065, A2 => n456, A3 => n454, A4 => n455, ZN
                           => n1059);
   U945 : AND4_X1 port map( A1 => n453, A2 => n452, A3 => n451, A4 => n450, ZN 
                           => n1065);
   U946 : AND4_X1 port map( A1 => n1066, A2 => n463, A3 => n461, A4 => n462, ZN
                           => n1058);
   U947 : AND4_X1 port map( A1 => n460, A2 => n459, A3 => n458, A4 => n457, ZN 
                           => n1066);
   U948 : OAI211_X1 port map( C1 => n1130, C2 => n877, A => n934, B => 
                           fill_port, ZN => n1056);
   U949 : INV_X1 port map( A => memory_response, ZN => n877);
   U950 : XOR2_X1 port map( A => n1067, B => n1068, Z => addr_r_4_port);
   U951 : XNOR2_X1 port map( A => address_w(4), B => n1069, ZN => n1068);
   U952 : OAI21_X1 port map( B1 => n1070, B2 => n1071, A => n1072, ZN => n1069)
                           ;
   U953 : OAI21_X1 port map( B1 => n1073, B2 => n1074, A => address_w(3), ZN =>
                           n1072);
   U954 : INV_X1 port map( A => n1073, ZN => n1071);
   U955 : NAND2_X1 port map( A1 => n1075, A2 => cwp_o_1_port, ZN => n1067);
   U956 : XOR2_X1 port map( A => n1076, B => n1074, Z => addr_r_3_port);
   U957 : INV_X1 port map( A => n1070, ZN => n1074);
   U958 : NAND2_X1 port map( A1 => n1077, A2 => n1078, ZN => n1070);
   U959 : XOR2_X1 port map( A => address_w(3), B => n1073, Z => n1076);
   U960 : OAI21_X1 port map( B1 => n1079, B2 => n1080, A => n1081, ZN => n1073)
                           ;
   U961 : OAI21_X1 port map( B1 => n1082, B2 => n1083, A => address_w(2), ZN =>
                           n1081);
   U962 : INV_X1 port map( A => n1079, ZN => n1083);
   U963 : INV_X1 port map( A => n1080, ZN => n1082);
   U964 : XOR2_X1 port map( A => n1079, B => n1084, Z => addr_r_2_port);
   U965 : XOR2_X1 port map( A => n1080, B => address_w(2), Z => n1084);
   U966 : NAND2_X1 port map( A1 => address_w(1), A2 => n1075, ZN => n1080);
   U967 : NAND2_X1 port map( A1 => n1085, A2 => n1078, ZN => n1079);
   U968 : XOR2_X1 port map( A => address_w(1), B => n1075, Z => addr_r_1_port);
   U969 : AND2_X1 port map( A1 => N1274, A2 => n1078, ZN => n1075);
   U970 : OR2_X1 port map( A1 => address_w(3), A2 => address_w(4), ZN => n1078)
                           ;
   U971 : XOR2_X1 port map( A => n1086, B => n1087, Z => addr_2_4_port);
   U972 : XNOR2_X1 port map( A => address_r_2(4), B => n1088, ZN => n1087);
   U973 : OAI21_X1 port map( B1 => n1089, B2 => n1090, A => n1091, ZN => n1088)
                           ;
   U974 : OAI21_X1 port map( B1 => n1092, B2 => n1093, A => address_r_2(3), ZN 
                           => n1091);
   U975 : INV_X1 port map( A => n1092, ZN => n1090);
   U976 : NAND2_X1 port map( A1 => n1094, A2 => cwp_o_1_port, ZN => n1086);
   U977 : XOR2_X1 port map( A => n1095, B => n1093, Z => addr_2_3_port);
   U978 : INV_X1 port map( A => n1089, ZN => n1093);
   U979 : NAND2_X1 port map( A1 => n1077, A2 => n1096, ZN => n1089);
   U980 : XOR2_X1 port map( A => address_r_2(3), B => n1092, Z => n1095);
   U981 : OAI21_X1 port map( B1 => n1097, B2 => n1098, A => n1099, ZN => n1092)
                           ;
   U982 : OAI21_X1 port map( B1 => n1100, B2 => n1101, A => address_r_2(2), ZN 
                           => n1099);
   U983 : INV_X1 port map( A => n1097, ZN => n1101);
   U984 : INV_X1 port map( A => n1098, ZN => n1100);
   U985 : XOR2_X1 port map( A => n1097, B => n1102, Z => addr_2_2_port);
   U986 : XOR2_X1 port map( A => n1098, B => address_r_2(2), Z => n1102);
   U987 : NAND2_X1 port map( A1 => address_r_2(1), A2 => n1094, ZN => n1098);
   U988 : NAND2_X1 port map( A1 => n1085, A2 => n1096, ZN => n1097);
   U989 : XOR2_X1 port map( A => address_r_2(1), B => n1094, Z => addr_2_1_port
                           );
   U990 : AND2_X1 port map( A1 => N1274, A2 => n1096, ZN => n1094);
   U991 : OR2_X1 port map( A1 => address_r_2(3), A2 => address_r_2(4), ZN => 
                           n1096);
   U992 : XOR2_X1 port map( A => n1103, B => n1104, Z => addr_1_4_port);
   U993 : XNOR2_X1 port map( A => address_r_1(4), B => n1105, ZN => n1104);
   U994 : OAI21_X1 port map( B1 => n1106, B2 => n1107, A => n1108, ZN => n1105)
                           ;
   U995 : OAI21_X1 port map( B1 => n1109, B2 => n1110, A => address_r_1(3), ZN 
                           => n1108);
   U996 : INV_X1 port map( A => n1109, ZN => n1107);
   U997 : NAND2_X1 port map( A1 => n1111, A2 => cwp_o_1_port, ZN => n1103);
   U998 : XOR2_X1 port map( A => n1112, B => n1110, Z => addr_1_3_port);
   U999 : INV_X1 port map( A => n1106, ZN => n1110);
   U1000 : NAND2_X1 port map( A1 => n1077, A2 => n1113, ZN => n1106);
   U1001 : XOR2_X1 port map( A => address_r_1(3), B => n1109, Z => n1112);
   U1002 : OAI21_X1 port map( B1 => n1114, B2 => n1115, A => n1116, ZN => n1109
                           );
   U1003 : OAI21_X1 port map( B1 => n1117, B2 => n1118, A => address_r_1(2), ZN
                           => n1116);
   U1004 : INV_X1 port map( A => n1114, ZN => n1118);
   U1005 : INV_X1 port map( A => n1115, ZN => n1117);
   U1006 : XOR2_X1 port map( A => n1114, B => n1119, Z => addr_1_2_port);
   U1007 : XOR2_X1 port map( A => n1115, B => address_r_1(2), Z => n1119);
   U1008 : NAND2_X1 port map( A1 => address_r_1(1), A2 => n1111, ZN => n1115);
   U1009 : NAND2_X1 port map( A1 => n1085, A2 => n1113, ZN => n1114);
   U1010 : INV_X1 port map( A => n1120, ZN => n1085);
   U1011 : AOI21_X1 port map( B1 => N1274, B2 => n273_port, A => n1077, ZN => 
                           n1120);
   U1012 : NOR2_X1 port map( A1 => N1274, A2 => n273_port, ZN => n1077);
   U1013 : XOR2_X1 port map( A => address_r_1(1), B => n1111, Z => 
                           addr_1_1_port);
   U1014 : AND2_X1 port map( A1 => N1274, A2 => n1113, ZN => n1111);
   U1015 : OR2_X1 port map( A1 => address_r_1(3), A2 => address_r_1(4), ZN => 
                           n1113);
   U1016 : MUX2_X1 port map( A => n1053, B => ret, S => n1052, Z => U3_U6_Z_0);
   U1017 : INV_X1 port map( A => call, ZN => n1052);
   U1018 : AND4_X1 port map( A1 => n431, A2 => n966, A3 => n466, A4 => n432, ZN
                           => n1053);
   U1019 : AND4_X1 port map( A1 => n1121, A2 => n1122, A3 => n1123, A4 => n1124
                           , ZN => n966);
   U1020 : NOR2_X1 port map( A1 => n1125, A2 => n1126, ZN => n1124);
   U1021 : NAND4_X1 port map( A1 => n409, A2 => n408, A3 => n407, A4 => n406, 
                           ZN => n1126);
   U1022 : NAND4_X1 port map( A1 => n405, A2 => n404, A3 => n403, A4 => n402, 
                           ZN => n1125);
   U1023 : AND4_X1 port map( A1 => n1127, A2 => n416, A3 => n414, A4 => n415, 
                           ZN => n1123);
   U1024 : AND4_X1 port map( A1 => n413, A2 => n412, A3 => n411, A4 => n410, ZN
                           => n1127);
   U1025 : AND4_X1 port map( A1 => n1128, A2 => n423, A3 => n421, A4 => n422, 
                           ZN => n1122);
   U1026 : AND4_X1 port map( A1 => n420, A2 => n419, A3 => n418, A4 => n417, ZN
                           => n1128);
   U1027 : AND4_X1 port map( A1 => n1129, A2 => n430, A3 => n428, A4 => n429, 
                           ZN => n1121);
   U1028 : AND4_X1 port map( A1 => n427, A2 => n426, A3 => n425, A4 => n424, ZN
                           => n1129);
   U1029 : INV_X1 port map( A => n934, ZN => N1006);
   U1030 : AOI21_X1 port map( B1 => n1044, B2 => n926, A => rest, ZN => n934);
   U1031 : NAND2_X1 port map( A1 => n1131, A2 => n1132, ZN => n926);
   U1032 : INV_X1 port map( A => n879, ZN => n1044);
   U1033 : NOR3_X1 port map( A1 => n1132, A2 => n1131, A3 => n799, ZN => n879);

end SYN_Behavioral;
