
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file.all;

entity register_file is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file;

architecture SYN_A of register_file is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal REGISTERS_0_63_port, REGISTERS_0_62_port, REGISTERS_0_61_port, 
      REGISTERS_0_60_port, REGISTERS_0_59_port, REGISTERS_0_58_port, 
      REGISTERS_0_57_port, REGISTERS_0_56_port, REGISTERS_0_55_port, 
      REGISTERS_0_54_port, REGISTERS_0_53_port, REGISTERS_0_52_port, 
      REGISTERS_0_51_port, REGISTERS_0_50_port, REGISTERS_0_49_port, 
      REGISTERS_0_48_port, REGISTERS_0_47_port, REGISTERS_0_46_port, 
      REGISTERS_0_45_port, REGISTERS_0_44_port, REGISTERS_0_43_port, 
      REGISTERS_0_42_port, REGISTERS_0_41_port, REGISTERS_0_40_port, 
      REGISTERS_0_39_port, REGISTERS_0_38_port, REGISTERS_0_37_port, 
      REGISTERS_0_36_port, REGISTERS_0_35_port, REGISTERS_0_34_port, 
      REGISTERS_0_33_port, REGISTERS_0_32_port, REGISTERS_0_31_port, 
      REGISTERS_0_30_port, REGISTERS_0_29_port, REGISTERS_0_28_port, 
      REGISTERS_0_27_port, REGISTERS_0_26_port, REGISTERS_0_25_port, 
      REGISTERS_0_24_port, REGISTERS_0_23_port, REGISTERS_0_22_port, 
      REGISTERS_0_21_port, REGISTERS_0_20_port, REGISTERS_0_19_port, 
      REGISTERS_0_18_port, REGISTERS_0_17_port, REGISTERS_0_16_port, 
      REGISTERS_0_15_port, REGISTERS_0_14_port, REGISTERS_0_13_port, 
      REGISTERS_0_12_port, REGISTERS_0_11_port, REGISTERS_0_10_port, 
      REGISTERS_0_9_port, REGISTERS_0_8_port, REGISTERS_0_7_port, 
      REGISTERS_0_6_port, REGISTERS_0_5_port, REGISTERS_0_4_port, 
      REGISTERS_0_3_port, REGISTERS_0_2_port, REGISTERS_0_1_port, 
      REGISTERS_0_0_port, REGISTERS_1_63_port, REGISTERS_1_62_port, 
      REGISTERS_1_61_port, REGISTERS_1_60_port, REGISTERS_1_59_port, 
      REGISTERS_1_58_port, REGISTERS_1_57_port, REGISTERS_1_56_port, 
      REGISTERS_1_55_port, REGISTERS_1_54_port, REGISTERS_1_53_port, 
      REGISTERS_1_52_port, REGISTERS_1_51_port, REGISTERS_1_50_port, 
      REGISTERS_1_49_port, REGISTERS_1_48_port, REGISTERS_1_47_port, 
      REGISTERS_1_46_port, REGISTERS_1_45_port, REGISTERS_1_44_port, 
      REGISTERS_1_43_port, REGISTERS_1_42_port, REGISTERS_1_41_port, 
      REGISTERS_1_40_port, REGISTERS_1_39_port, REGISTERS_1_38_port, 
      REGISTERS_1_37_port, REGISTERS_1_36_port, REGISTERS_1_35_port, 
      REGISTERS_1_34_port, REGISTERS_1_33_port, REGISTERS_1_32_port, 
      REGISTERS_1_31_port, REGISTERS_1_30_port, REGISTERS_1_29_port, 
      REGISTERS_1_28_port, REGISTERS_1_27_port, REGISTERS_1_26_port, 
      REGISTERS_1_25_port, REGISTERS_1_24_port, REGISTERS_1_23_port, 
      REGISTERS_1_22_port, REGISTERS_1_21_port, REGISTERS_1_20_port, 
      REGISTERS_1_19_port, REGISTERS_1_18_port, REGISTERS_1_17_port, 
      REGISTERS_1_16_port, REGISTERS_1_15_port, REGISTERS_1_14_port, 
      REGISTERS_1_13_port, REGISTERS_1_12_port, REGISTERS_1_11_port, 
      REGISTERS_1_10_port, REGISTERS_1_9_port, REGISTERS_1_8_port, 
      REGISTERS_1_7_port, REGISTERS_1_6_port, REGISTERS_1_5_port, 
      REGISTERS_1_4_port, REGISTERS_1_3_port, REGISTERS_1_2_port, 
      REGISTERS_1_1_port, REGISTERS_1_0_port, REGISTERS_2_63_port, 
      REGISTERS_2_62_port, REGISTERS_2_61_port, REGISTERS_2_60_port, 
      REGISTERS_2_59_port, REGISTERS_2_58_port, REGISTERS_2_57_port, 
      REGISTERS_2_56_port, REGISTERS_2_55_port, REGISTERS_2_54_port, 
      REGISTERS_2_53_port, REGISTERS_2_52_port, REGISTERS_2_51_port, 
      REGISTERS_2_50_port, REGISTERS_2_49_port, REGISTERS_2_48_port, 
      REGISTERS_2_47_port, REGISTERS_2_46_port, REGISTERS_2_45_port, 
      REGISTERS_2_44_port, REGISTERS_2_43_port, REGISTERS_2_42_port, 
      REGISTERS_2_41_port, REGISTERS_2_40_port, REGISTERS_2_39_port, 
      REGISTERS_2_38_port, REGISTERS_2_37_port, REGISTERS_2_36_port, 
      REGISTERS_2_35_port, REGISTERS_2_34_port, REGISTERS_2_33_port, 
      REGISTERS_2_32_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_63_port, REGISTERS_3_62_port, REGISTERS_3_61_port, 
      REGISTERS_3_60_port, REGISTERS_3_59_port, REGISTERS_3_58_port, 
      REGISTERS_3_57_port, REGISTERS_3_56_port, REGISTERS_3_55_port, 
      REGISTERS_3_54_port, REGISTERS_3_53_port, REGISTERS_3_52_port, 
      REGISTERS_3_51_port, REGISTERS_3_50_port, REGISTERS_3_49_port, 
      REGISTERS_3_48_port, REGISTERS_3_47_port, REGISTERS_3_46_port, 
      REGISTERS_3_45_port, REGISTERS_3_44_port, REGISTERS_3_43_port, 
      REGISTERS_3_42_port, REGISTERS_3_41_port, REGISTERS_3_40_port, 
      REGISTERS_3_39_port, REGISTERS_3_38_port, REGISTERS_3_37_port, 
      REGISTERS_3_36_port, REGISTERS_3_35_port, REGISTERS_3_34_port, 
      REGISTERS_3_33_port, REGISTERS_3_32_port, REGISTERS_3_31_port, 
      REGISTERS_3_30_port, REGISTERS_3_29_port, REGISTERS_3_28_port, 
      REGISTERS_3_27_port, REGISTERS_3_26_port, REGISTERS_3_25_port, 
      REGISTERS_3_24_port, REGISTERS_3_23_port, REGISTERS_3_22_port, 
      REGISTERS_3_21_port, REGISTERS_3_20_port, REGISTERS_3_19_port, 
      REGISTERS_3_18_port, REGISTERS_3_17_port, REGISTERS_3_16_port, 
      REGISTERS_3_15_port, REGISTERS_3_14_port, REGISTERS_3_13_port, 
      REGISTERS_3_12_port, REGISTERS_3_11_port, REGISTERS_3_10_port, 
      REGISTERS_3_9_port, REGISTERS_3_8_port, REGISTERS_3_7_port, 
      REGISTERS_3_6_port, REGISTERS_3_5_port, REGISTERS_3_4_port, 
      REGISTERS_3_3_port, REGISTERS_3_2_port, REGISTERS_3_1_port, 
      REGISTERS_3_0_port, REGISTERS_4_63_port, REGISTERS_4_62_port, 
      REGISTERS_4_61_port, REGISTERS_4_60_port, REGISTERS_4_59_port, 
      REGISTERS_4_58_port, REGISTERS_4_57_port, REGISTERS_4_56_port, 
      REGISTERS_4_55_port, REGISTERS_4_54_port, REGISTERS_4_53_port, 
      REGISTERS_4_52_port, REGISTERS_4_51_port, REGISTERS_4_50_port, 
      REGISTERS_4_49_port, REGISTERS_4_48_port, REGISTERS_4_47_port, 
      REGISTERS_4_46_port, REGISTERS_4_45_port, REGISTERS_4_44_port, 
      REGISTERS_4_43_port, REGISTERS_4_42_port, REGISTERS_4_41_port, 
      REGISTERS_4_40_port, REGISTERS_4_39_port, REGISTERS_4_38_port, 
      REGISTERS_4_37_port, REGISTERS_4_36_port, REGISTERS_4_35_port, 
      REGISTERS_4_34_port, REGISTERS_4_33_port, REGISTERS_4_32_port, 
      REGISTERS_4_31_port, REGISTERS_4_30_port, REGISTERS_4_29_port, 
      REGISTERS_4_28_port, REGISTERS_4_27_port, REGISTERS_4_26_port, 
      REGISTERS_4_25_port, REGISTERS_4_24_port, REGISTERS_4_23_port, 
      REGISTERS_4_22_port, REGISTERS_4_21_port, REGISTERS_4_20_port, 
      REGISTERS_4_19_port, REGISTERS_4_18_port, REGISTERS_4_17_port, 
      REGISTERS_4_16_port, REGISTERS_4_15_port, REGISTERS_4_14_port, 
      REGISTERS_4_13_port, REGISTERS_4_12_port, REGISTERS_4_11_port, 
      REGISTERS_4_10_port, REGISTERS_4_9_port, REGISTERS_4_8_port, 
      REGISTERS_4_7_port, REGISTERS_4_6_port, REGISTERS_4_5_port, 
      REGISTERS_4_4_port, REGISTERS_4_3_port, REGISTERS_4_2_port, 
      REGISTERS_4_1_port, REGISTERS_4_0_port, REGISTERS_5_63_port, 
      REGISTERS_5_62_port, REGISTERS_5_61_port, REGISTERS_5_60_port, 
      REGISTERS_5_59_port, REGISTERS_5_58_port, REGISTERS_5_57_port, 
      REGISTERS_5_56_port, REGISTERS_5_55_port, REGISTERS_5_54_port, 
      REGISTERS_5_53_port, REGISTERS_5_52_port, REGISTERS_5_51_port, 
      REGISTERS_5_50_port, REGISTERS_5_49_port, REGISTERS_5_48_port, 
      REGISTERS_5_47_port, REGISTERS_5_46_port, REGISTERS_5_45_port, 
      REGISTERS_5_44_port, REGISTERS_5_43_port, REGISTERS_5_42_port, 
      REGISTERS_5_41_port, REGISTERS_5_40_port, REGISTERS_5_39_port, 
      REGISTERS_5_38_port, REGISTERS_5_37_port, REGISTERS_5_36_port, 
      REGISTERS_5_35_port, REGISTERS_5_34_port, REGISTERS_5_33_port, 
      REGISTERS_5_32_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_63_port, REGISTERS_6_62_port, REGISTERS_6_61_port, 
      REGISTERS_6_60_port, REGISTERS_6_59_port, REGISTERS_6_58_port, 
      REGISTERS_6_57_port, REGISTERS_6_56_port, REGISTERS_6_55_port, 
      REGISTERS_6_54_port, REGISTERS_6_53_port, REGISTERS_6_52_port, 
      REGISTERS_6_51_port, REGISTERS_6_50_port, REGISTERS_6_49_port, 
      REGISTERS_6_48_port, REGISTERS_6_47_port, REGISTERS_6_46_port, 
      REGISTERS_6_45_port, REGISTERS_6_44_port, REGISTERS_6_43_port, 
      REGISTERS_6_42_port, REGISTERS_6_41_port, REGISTERS_6_40_port, 
      REGISTERS_6_39_port, REGISTERS_6_38_port, REGISTERS_6_37_port, 
      REGISTERS_6_36_port, REGISTERS_6_35_port, REGISTERS_6_34_port, 
      REGISTERS_6_33_port, REGISTERS_6_32_port, REGISTERS_6_31_port, 
      REGISTERS_6_30_port, REGISTERS_6_29_port, REGISTERS_6_28_port, 
      REGISTERS_6_27_port, REGISTERS_6_26_port, REGISTERS_6_25_port, 
      REGISTERS_6_24_port, REGISTERS_6_23_port, REGISTERS_6_22_port, 
      REGISTERS_6_21_port, REGISTERS_6_20_port, REGISTERS_6_19_port, 
      REGISTERS_6_18_port, REGISTERS_6_17_port, REGISTERS_6_16_port, 
      REGISTERS_6_15_port, REGISTERS_6_14_port, REGISTERS_6_13_port, 
      REGISTERS_6_12_port, REGISTERS_6_11_port, REGISTERS_6_10_port, 
      REGISTERS_6_9_port, REGISTERS_6_8_port, REGISTERS_6_7_port, 
      REGISTERS_6_6_port, REGISTERS_6_5_port, REGISTERS_6_4_port, 
      REGISTERS_6_3_port, REGISTERS_6_2_port, REGISTERS_6_1_port, 
      REGISTERS_6_0_port, REGISTERS_7_63_port, REGISTERS_7_62_port, 
      REGISTERS_7_61_port, REGISTERS_7_60_port, REGISTERS_7_59_port, 
      REGISTERS_7_58_port, REGISTERS_7_57_port, REGISTERS_7_56_port, 
      REGISTERS_7_55_port, REGISTERS_7_54_port, REGISTERS_7_53_port, 
      REGISTERS_7_52_port, REGISTERS_7_51_port, REGISTERS_7_50_port, 
      REGISTERS_7_49_port, REGISTERS_7_48_port, REGISTERS_7_47_port, 
      REGISTERS_7_46_port, REGISTERS_7_45_port, REGISTERS_7_44_port, 
      REGISTERS_7_43_port, REGISTERS_7_42_port, REGISTERS_7_41_port, 
      REGISTERS_7_40_port, REGISTERS_7_39_port, REGISTERS_7_38_port, 
      REGISTERS_7_37_port, REGISTERS_7_36_port, REGISTERS_7_35_port, 
      REGISTERS_7_34_port, REGISTERS_7_33_port, REGISTERS_7_32_port, 
      REGISTERS_7_31_port, REGISTERS_7_30_port, REGISTERS_7_29_port, 
      REGISTERS_7_28_port, REGISTERS_7_27_port, REGISTERS_7_26_port, 
      REGISTERS_7_25_port, REGISTERS_7_24_port, REGISTERS_7_23_port, 
      REGISTERS_7_22_port, REGISTERS_7_21_port, REGISTERS_7_20_port, 
      REGISTERS_7_19_port, REGISTERS_7_18_port, REGISTERS_7_17_port, 
      REGISTERS_7_16_port, REGISTERS_7_15_port, REGISTERS_7_14_port, 
      REGISTERS_7_13_port, REGISTERS_7_12_port, REGISTERS_7_11_port, 
      REGISTERS_7_10_port, REGISTERS_7_9_port, REGISTERS_7_8_port, 
      REGISTERS_7_7_port, REGISTERS_7_6_port, REGISTERS_7_5_port, 
      REGISTERS_7_4_port, REGISTERS_7_3_port, REGISTERS_7_2_port, 
      REGISTERS_7_1_port, REGISTERS_7_0_port, REGISTERS_8_63_port, 
      REGISTERS_8_62_port, REGISTERS_8_61_port, REGISTERS_8_60_port, 
      REGISTERS_8_59_port, REGISTERS_8_58_port, REGISTERS_8_57_port, 
      REGISTERS_8_56_port, REGISTERS_8_55_port, REGISTERS_8_54_port, 
      REGISTERS_8_53_port, REGISTERS_8_52_port, REGISTERS_8_51_port, 
      REGISTERS_8_50_port, REGISTERS_8_49_port, REGISTERS_8_48_port, 
      REGISTERS_8_47_port, REGISTERS_8_46_port, REGISTERS_8_45_port, 
      REGISTERS_8_44_port, REGISTERS_8_43_port, REGISTERS_8_42_port, 
      REGISTERS_8_41_port, REGISTERS_8_40_port, REGISTERS_8_39_port, 
      REGISTERS_8_38_port, REGISTERS_8_37_port, REGISTERS_8_36_port, 
      REGISTERS_8_35_port, REGISTERS_8_34_port, REGISTERS_8_33_port, 
      REGISTERS_8_32_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_63_port, REGISTERS_9_62_port, REGISTERS_9_61_port, 
      REGISTERS_9_60_port, REGISTERS_9_59_port, REGISTERS_9_58_port, 
      REGISTERS_9_57_port, REGISTERS_9_56_port, REGISTERS_9_55_port, 
      REGISTERS_9_54_port, REGISTERS_9_53_port, REGISTERS_9_52_port, 
      REGISTERS_9_51_port, REGISTERS_9_50_port, REGISTERS_9_49_port, 
      REGISTERS_9_48_port, REGISTERS_9_47_port, REGISTERS_9_46_port, 
      REGISTERS_9_45_port, REGISTERS_9_44_port, REGISTERS_9_43_port, 
      REGISTERS_9_42_port, REGISTERS_9_41_port, REGISTERS_9_40_port, 
      REGISTERS_9_39_port, REGISTERS_9_38_port, REGISTERS_9_37_port, 
      REGISTERS_9_36_port, REGISTERS_9_35_port, REGISTERS_9_34_port, 
      REGISTERS_9_33_port, REGISTERS_9_32_port, REGISTERS_9_31_port, 
      REGISTERS_9_30_port, REGISTERS_9_29_port, REGISTERS_9_28_port, 
      REGISTERS_9_27_port, REGISTERS_9_26_port, REGISTERS_9_25_port, 
      REGISTERS_9_24_port, REGISTERS_9_23_port, REGISTERS_9_22_port, 
      REGISTERS_9_21_port, REGISTERS_9_20_port, REGISTERS_9_19_port, 
      REGISTERS_9_18_port, REGISTERS_9_17_port, REGISTERS_9_16_port, 
      REGISTERS_9_15_port, REGISTERS_9_14_port, REGISTERS_9_13_port, 
      REGISTERS_9_12_port, REGISTERS_9_11_port, REGISTERS_9_10_port, 
      REGISTERS_9_9_port, REGISTERS_9_8_port, REGISTERS_9_7_port, 
      REGISTERS_9_6_port, REGISTERS_9_5_port, REGISTERS_9_4_port, 
      REGISTERS_9_3_port, REGISTERS_9_2_port, REGISTERS_9_1_port, 
      REGISTERS_9_0_port, REGISTERS_10_63_port, REGISTERS_10_62_port, 
      REGISTERS_10_61_port, REGISTERS_10_60_port, REGISTERS_10_59_port, 
      REGISTERS_10_58_port, REGISTERS_10_57_port, REGISTERS_10_56_port, 
      REGISTERS_10_55_port, REGISTERS_10_54_port, REGISTERS_10_53_port, 
      REGISTERS_10_52_port, REGISTERS_10_51_port, REGISTERS_10_50_port, 
      REGISTERS_10_49_port, REGISTERS_10_48_port, REGISTERS_10_47_port, 
      REGISTERS_10_46_port, REGISTERS_10_45_port, REGISTERS_10_44_port, 
      REGISTERS_10_43_port, REGISTERS_10_42_port, REGISTERS_10_41_port, 
      REGISTERS_10_40_port, REGISTERS_10_39_port, REGISTERS_10_38_port, 
      REGISTERS_10_37_port, REGISTERS_10_36_port, REGISTERS_10_35_port, 
      REGISTERS_10_34_port, REGISTERS_10_33_port, REGISTERS_10_32_port, 
      REGISTERS_10_31_port, REGISTERS_10_30_port, REGISTERS_10_29_port, 
      REGISTERS_10_28_port, REGISTERS_10_27_port, REGISTERS_10_26_port, 
      REGISTERS_10_25_port, REGISTERS_10_24_port, REGISTERS_10_23_port, 
      REGISTERS_10_22_port, REGISTERS_10_21_port, REGISTERS_10_20_port, 
      REGISTERS_10_19_port, REGISTERS_10_18_port, REGISTERS_10_17_port, 
      REGISTERS_10_16_port, REGISTERS_10_15_port, REGISTERS_10_14_port, 
      REGISTERS_10_13_port, REGISTERS_10_12_port, REGISTERS_10_11_port, 
      REGISTERS_10_10_port, REGISTERS_10_9_port, REGISTERS_10_8_port, 
      REGISTERS_10_7_port, REGISTERS_10_6_port, REGISTERS_10_5_port, 
      REGISTERS_10_4_port, REGISTERS_10_3_port, REGISTERS_10_2_port, 
      REGISTERS_10_1_port, REGISTERS_10_0_port, REGISTERS_11_63_port, 
      REGISTERS_11_62_port, REGISTERS_11_61_port, REGISTERS_11_60_port, 
      REGISTERS_11_59_port, REGISTERS_11_58_port, REGISTERS_11_57_port, 
      REGISTERS_11_56_port, REGISTERS_11_55_port, REGISTERS_11_54_port, 
      REGISTERS_11_53_port, REGISTERS_11_52_port, REGISTERS_11_51_port, 
      REGISTERS_11_50_port, REGISTERS_11_49_port, REGISTERS_11_48_port, 
      REGISTERS_11_47_port, REGISTERS_11_46_port, REGISTERS_11_45_port, 
      REGISTERS_11_44_port, REGISTERS_11_43_port, REGISTERS_11_42_port, 
      REGISTERS_11_41_port, REGISTERS_11_40_port, REGISTERS_11_39_port, 
      REGISTERS_11_38_port, REGISTERS_11_37_port, REGISTERS_11_36_port, 
      REGISTERS_11_35_port, REGISTERS_11_34_port, REGISTERS_11_33_port, 
      REGISTERS_11_32_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_63_port, REGISTERS_12_62_port, REGISTERS_12_61_port, 
      REGISTERS_12_60_port, REGISTERS_12_59_port, REGISTERS_12_58_port, 
      REGISTERS_12_57_port, REGISTERS_12_56_port, REGISTERS_12_55_port, 
      REGISTERS_12_54_port, REGISTERS_12_53_port, REGISTERS_12_52_port, 
      REGISTERS_12_51_port, REGISTERS_12_50_port, REGISTERS_12_49_port, 
      REGISTERS_12_48_port, REGISTERS_12_47_port, REGISTERS_12_46_port, 
      REGISTERS_12_45_port, REGISTERS_12_44_port, REGISTERS_12_43_port, 
      REGISTERS_12_42_port, REGISTERS_12_41_port, REGISTERS_12_40_port, 
      REGISTERS_12_39_port, REGISTERS_12_38_port, REGISTERS_12_37_port, 
      REGISTERS_12_36_port, REGISTERS_12_35_port, REGISTERS_12_34_port, 
      REGISTERS_12_33_port, REGISTERS_12_32_port, REGISTERS_12_31_port, 
      REGISTERS_12_30_port, REGISTERS_12_29_port, REGISTERS_12_28_port, 
      REGISTERS_12_27_port, REGISTERS_12_26_port, REGISTERS_12_25_port, 
      REGISTERS_12_24_port, REGISTERS_12_23_port, REGISTERS_12_22_port, 
      REGISTERS_12_21_port, REGISTERS_12_20_port, REGISTERS_12_19_port, 
      REGISTERS_12_18_port, REGISTERS_12_17_port, REGISTERS_12_16_port, 
      REGISTERS_12_15_port, REGISTERS_12_14_port, REGISTERS_12_13_port, 
      REGISTERS_12_12_port, REGISTERS_12_11_port, REGISTERS_12_10_port, 
      REGISTERS_12_9_port, REGISTERS_12_8_port, REGISTERS_12_7_port, 
      REGISTERS_12_6_port, REGISTERS_12_5_port, REGISTERS_12_4_port, 
      REGISTERS_12_3_port, REGISTERS_12_2_port, REGISTERS_12_1_port, 
      REGISTERS_12_0_port, REGISTERS_13_63_port, REGISTERS_13_62_port, 
      REGISTERS_13_61_port, REGISTERS_13_60_port, REGISTERS_13_59_port, 
      REGISTERS_13_58_port, REGISTERS_13_57_port, REGISTERS_13_56_port, 
      REGISTERS_13_55_port, REGISTERS_13_54_port, REGISTERS_13_53_port, 
      REGISTERS_13_52_port, REGISTERS_13_51_port, REGISTERS_13_50_port, 
      REGISTERS_13_49_port, REGISTERS_13_48_port, REGISTERS_13_47_port, 
      REGISTERS_13_46_port, REGISTERS_13_45_port, REGISTERS_13_44_port, 
      REGISTERS_13_43_port, REGISTERS_13_42_port, REGISTERS_13_41_port, 
      REGISTERS_13_40_port, REGISTERS_13_39_port, REGISTERS_13_38_port, 
      REGISTERS_13_37_port, REGISTERS_13_36_port, REGISTERS_13_35_port, 
      REGISTERS_13_34_port, REGISTERS_13_33_port, REGISTERS_13_32_port, 
      REGISTERS_13_31_port, REGISTERS_13_30_port, REGISTERS_13_29_port, 
      REGISTERS_13_28_port, REGISTERS_13_27_port, REGISTERS_13_26_port, 
      REGISTERS_13_25_port, REGISTERS_13_24_port, REGISTERS_13_23_port, 
      REGISTERS_13_22_port, REGISTERS_13_21_port, REGISTERS_13_20_port, 
      REGISTERS_13_19_port, REGISTERS_13_18_port, REGISTERS_13_17_port, 
      REGISTERS_13_16_port, REGISTERS_13_15_port, REGISTERS_13_14_port, 
      REGISTERS_13_13_port, REGISTERS_13_12_port, REGISTERS_13_11_port, 
      REGISTERS_13_10_port, REGISTERS_13_9_port, REGISTERS_13_8_port, 
      REGISTERS_13_7_port, REGISTERS_13_6_port, REGISTERS_13_5_port, 
      REGISTERS_13_4_port, REGISTERS_13_3_port, REGISTERS_13_2_port, 
      REGISTERS_13_1_port, REGISTERS_13_0_port, REGISTERS_14_63_port, 
      REGISTERS_14_62_port, REGISTERS_14_61_port, REGISTERS_14_60_port, 
      REGISTERS_14_59_port, REGISTERS_14_58_port, REGISTERS_14_57_port, 
      REGISTERS_14_56_port, REGISTERS_14_55_port, REGISTERS_14_54_port, 
      REGISTERS_14_53_port, REGISTERS_14_52_port, REGISTERS_14_51_port, 
      REGISTERS_14_50_port, REGISTERS_14_49_port, REGISTERS_14_48_port, 
      REGISTERS_14_47_port, REGISTERS_14_46_port, REGISTERS_14_45_port, 
      REGISTERS_14_44_port, REGISTERS_14_43_port, REGISTERS_14_42_port, 
      REGISTERS_14_41_port, REGISTERS_14_40_port, REGISTERS_14_39_port, 
      REGISTERS_14_38_port, REGISTERS_14_37_port, REGISTERS_14_36_port, 
      REGISTERS_14_35_port, REGISTERS_14_34_port, REGISTERS_14_33_port, 
      REGISTERS_14_32_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_63_port, REGISTERS_15_62_port, REGISTERS_15_61_port, 
      REGISTERS_15_60_port, REGISTERS_15_59_port, REGISTERS_15_58_port, 
      REGISTERS_15_57_port, REGISTERS_15_56_port, REGISTERS_15_55_port, 
      REGISTERS_15_54_port, REGISTERS_15_53_port, REGISTERS_15_52_port, 
      REGISTERS_15_51_port, REGISTERS_15_50_port, REGISTERS_15_49_port, 
      REGISTERS_15_48_port, REGISTERS_15_47_port, REGISTERS_15_46_port, 
      REGISTERS_15_45_port, REGISTERS_15_44_port, REGISTERS_15_43_port, 
      REGISTERS_15_42_port, REGISTERS_15_41_port, REGISTERS_15_40_port, 
      REGISTERS_15_39_port, REGISTERS_15_38_port, REGISTERS_15_37_port, 
      REGISTERS_15_36_port, REGISTERS_15_35_port, REGISTERS_15_34_port, 
      REGISTERS_15_33_port, REGISTERS_15_32_port, REGISTERS_15_31_port, 
      REGISTERS_15_30_port, REGISTERS_15_29_port, REGISTERS_15_28_port, 
      REGISTERS_15_27_port, REGISTERS_15_26_port, REGISTERS_15_25_port, 
      REGISTERS_15_24_port, REGISTERS_15_23_port, REGISTERS_15_22_port, 
      REGISTERS_15_21_port, REGISTERS_15_20_port, REGISTERS_15_19_port, 
      REGISTERS_15_18_port, REGISTERS_15_17_port, REGISTERS_15_16_port, 
      REGISTERS_15_15_port, REGISTERS_15_14_port, REGISTERS_15_13_port, 
      REGISTERS_15_12_port, REGISTERS_15_11_port, REGISTERS_15_10_port, 
      REGISTERS_15_9_port, REGISTERS_15_8_port, REGISTERS_15_7_port, 
      REGISTERS_15_6_port, REGISTERS_15_5_port, REGISTERS_15_4_port, 
      REGISTERS_15_3_port, REGISTERS_15_2_port, REGISTERS_15_1_port, 
      REGISTERS_15_0_port, REGISTERS_16_63_port, REGISTERS_16_62_port, 
      REGISTERS_16_61_port, REGISTERS_16_60_port, REGISTERS_16_59_port, 
      REGISTERS_16_58_port, REGISTERS_16_57_port, REGISTERS_16_56_port, 
      REGISTERS_16_55_port, REGISTERS_16_54_port, REGISTERS_16_53_port, 
      REGISTERS_16_52_port, REGISTERS_16_51_port, REGISTERS_16_50_port, 
      REGISTERS_16_49_port, REGISTERS_16_48_port, REGISTERS_16_47_port, 
      REGISTERS_16_46_port, REGISTERS_16_45_port, REGISTERS_16_44_port, 
      REGISTERS_16_43_port, REGISTERS_16_42_port, REGISTERS_16_41_port, 
      REGISTERS_16_40_port, REGISTERS_16_39_port, REGISTERS_16_38_port, 
      REGISTERS_16_37_port, REGISTERS_16_36_port, REGISTERS_16_35_port, 
      REGISTERS_16_34_port, REGISTERS_16_33_port, REGISTERS_16_32_port, 
      REGISTERS_16_31_port, REGISTERS_16_30_port, REGISTERS_16_29_port, 
      REGISTERS_16_28_port, REGISTERS_16_27_port, REGISTERS_16_26_port, 
      REGISTERS_16_25_port, REGISTERS_16_24_port, REGISTERS_16_23_port, 
      REGISTERS_16_22_port, REGISTERS_16_21_port, REGISTERS_16_20_port, 
      REGISTERS_16_19_port, REGISTERS_16_18_port, REGISTERS_16_17_port, 
      REGISTERS_16_16_port, REGISTERS_16_15_port, REGISTERS_16_14_port, 
      REGISTERS_16_13_port, REGISTERS_16_12_port, REGISTERS_16_11_port, 
      REGISTERS_16_10_port, REGISTERS_16_9_port, REGISTERS_16_8_port, 
      REGISTERS_16_7_port, REGISTERS_16_6_port, REGISTERS_16_5_port, 
      REGISTERS_16_4_port, REGISTERS_16_3_port, REGISTERS_16_2_port, 
      REGISTERS_16_1_port, REGISTERS_16_0_port, REGISTERS_17_63_port, 
      REGISTERS_17_62_port, REGISTERS_17_61_port, REGISTERS_17_60_port, 
      REGISTERS_17_59_port, REGISTERS_17_58_port, REGISTERS_17_57_port, 
      REGISTERS_17_56_port, REGISTERS_17_55_port, REGISTERS_17_54_port, 
      REGISTERS_17_53_port, REGISTERS_17_52_port, REGISTERS_17_51_port, 
      REGISTERS_17_50_port, REGISTERS_17_49_port, REGISTERS_17_48_port, 
      REGISTERS_17_47_port, REGISTERS_17_46_port, REGISTERS_17_45_port, 
      REGISTERS_17_44_port, REGISTERS_17_43_port, REGISTERS_17_42_port, 
      REGISTERS_17_41_port, REGISTERS_17_40_port, REGISTERS_17_39_port, 
      REGISTERS_17_38_port, REGISTERS_17_37_port, REGISTERS_17_36_port, 
      REGISTERS_17_35_port, REGISTERS_17_34_port, REGISTERS_17_33_port, 
      REGISTERS_17_32_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_63_port, REGISTERS_18_62_port, REGISTERS_18_61_port, 
      REGISTERS_18_60_port, REGISTERS_18_59_port, REGISTERS_18_58_port, 
      REGISTERS_18_57_port, REGISTERS_18_56_port, REGISTERS_18_55_port, 
      REGISTERS_18_54_port, REGISTERS_18_53_port, REGISTERS_18_52_port, 
      REGISTERS_18_51_port, REGISTERS_18_50_port, REGISTERS_18_49_port, 
      REGISTERS_18_48_port, REGISTERS_18_47_port, REGISTERS_18_46_port, 
      REGISTERS_18_45_port, REGISTERS_18_44_port, REGISTERS_18_43_port, 
      REGISTERS_18_42_port, REGISTERS_18_41_port, REGISTERS_18_40_port, 
      REGISTERS_18_39_port, REGISTERS_18_38_port, REGISTERS_18_37_port, 
      REGISTERS_18_36_port, REGISTERS_18_35_port, REGISTERS_18_34_port, 
      REGISTERS_18_33_port, REGISTERS_18_32_port, REGISTERS_18_31_port, 
      REGISTERS_18_30_port, REGISTERS_18_29_port, REGISTERS_18_28_port, 
      REGISTERS_18_27_port, REGISTERS_18_26_port, REGISTERS_18_25_port, 
      REGISTERS_18_24_port, REGISTERS_18_23_port, REGISTERS_18_22_port, 
      REGISTERS_18_21_port, REGISTERS_18_20_port, REGISTERS_18_19_port, 
      REGISTERS_18_18_port, REGISTERS_18_17_port, REGISTERS_18_16_port, 
      REGISTERS_18_15_port, REGISTERS_18_14_port, REGISTERS_18_13_port, 
      REGISTERS_18_12_port, REGISTERS_18_11_port, REGISTERS_18_10_port, 
      REGISTERS_18_9_port, REGISTERS_18_8_port, REGISTERS_18_7_port, 
      REGISTERS_18_6_port, REGISTERS_18_5_port, REGISTERS_18_4_port, 
      REGISTERS_18_3_port, REGISTERS_18_2_port, REGISTERS_18_1_port, 
      REGISTERS_18_0_port, REGISTERS_19_63_port, REGISTERS_19_62_port, 
      REGISTERS_19_61_port, REGISTERS_19_60_port, REGISTERS_19_59_port, 
      REGISTERS_19_58_port, REGISTERS_19_57_port, REGISTERS_19_56_port, 
      REGISTERS_19_55_port, REGISTERS_19_54_port, REGISTERS_19_53_port, 
      REGISTERS_19_52_port, REGISTERS_19_51_port, REGISTERS_19_50_port, 
      REGISTERS_19_49_port, REGISTERS_19_48_port, REGISTERS_19_47_port, 
      REGISTERS_19_46_port, REGISTERS_19_45_port, REGISTERS_19_44_port, 
      REGISTERS_19_43_port, REGISTERS_19_42_port, REGISTERS_19_41_port, 
      REGISTERS_19_40_port, REGISTERS_19_39_port, REGISTERS_19_38_port, 
      REGISTERS_19_37_port, REGISTERS_19_36_port, REGISTERS_19_35_port, 
      REGISTERS_19_34_port, REGISTERS_19_33_port, REGISTERS_19_32_port, 
      REGISTERS_19_31_port, REGISTERS_19_30_port, REGISTERS_19_29_port, 
      REGISTERS_19_28_port, REGISTERS_19_27_port, REGISTERS_19_26_port, 
      REGISTERS_19_25_port, REGISTERS_19_24_port, REGISTERS_19_23_port, 
      REGISTERS_19_22_port, REGISTERS_19_21_port, REGISTERS_19_20_port, 
      REGISTERS_19_19_port, REGISTERS_19_18_port, REGISTERS_19_17_port, 
      REGISTERS_19_16_port, REGISTERS_19_15_port, REGISTERS_19_14_port, 
      REGISTERS_19_13_port, REGISTERS_19_12_port, REGISTERS_19_11_port, 
      REGISTERS_19_10_port, REGISTERS_19_9_port, REGISTERS_19_8_port, 
      REGISTERS_19_7_port, REGISTERS_19_6_port, REGISTERS_19_5_port, 
      REGISTERS_19_4_port, REGISTERS_19_3_port, REGISTERS_19_2_port, 
      REGISTERS_19_1_port, REGISTERS_19_0_port, REGISTERS_20_63_port, 
      REGISTERS_20_62_port, REGISTERS_20_61_port, REGISTERS_20_60_port, 
      REGISTERS_20_59_port, REGISTERS_20_58_port, REGISTERS_20_57_port, 
      REGISTERS_20_56_port, REGISTERS_20_55_port, REGISTERS_20_54_port, 
      REGISTERS_20_53_port, REGISTERS_20_52_port, REGISTERS_20_51_port, 
      REGISTERS_20_50_port, REGISTERS_20_49_port, REGISTERS_20_48_port, 
      REGISTERS_20_47_port, REGISTERS_20_46_port, REGISTERS_20_45_port, 
      REGISTERS_20_44_port, REGISTERS_20_43_port, REGISTERS_20_42_port, 
      REGISTERS_20_41_port, REGISTERS_20_40_port, REGISTERS_20_39_port, 
      REGISTERS_20_38_port, REGISTERS_20_37_port, REGISTERS_20_36_port, 
      REGISTERS_20_35_port, REGISTERS_20_34_port, REGISTERS_20_33_port, 
      REGISTERS_20_32_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_63_port, REGISTERS_21_62_port, REGISTERS_21_61_port, 
      REGISTERS_21_60_port, REGISTERS_21_59_port, REGISTERS_21_58_port, 
      REGISTERS_21_57_port, REGISTERS_21_56_port, REGISTERS_21_55_port, 
      REGISTERS_21_54_port, REGISTERS_21_53_port, REGISTERS_21_52_port, 
      REGISTERS_21_51_port, REGISTERS_21_50_port, REGISTERS_21_49_port, 
      REGISTERS_21_48_port, REGISTERS_21_47_port, REGISTERS_21_46_port, 
      REGISTERS_21_45_port, REGISTERS_21_44_port, REGISTERS_21_43_port, 
      REGISTERS_21_42_port, REGISTERS_21_41_port, REGISTERS_21_40_port, 
      REGISTERS_21_39_port, REGISTERS_21_38_port, REGISTERS_21_37_port, 
      REGISTERS_21_36_port, REGISTERS_21_35_port, REGISTERS_21_34_port, 
      REGISTERS_21_33_port, REGISTERS_21_32_port, REGISTERS_21_31_port, 
      REGISTERS_21_30_port, REGISTERS_21_29_port, REGISTERS_21_28_port, 
      REGISTERS_21_27_port, REGISTERS_21_26_port, REGISTERS_21_25_port, 
      REGISTERS_21_24_port, REGISTERS_21_23_port, REGISTERS_21_22_port, 
      REGISTERS_21_21_port, REGISTERS_21_20_port, REGISTERS_21_19_port, 
      REGISTERS_21_18_port, REGISTERS_21_17_port, REGISTERS_21_16_port, 
      REGISTERS_21_15_port, REGISTERS_21_14_port, REGISTERS_21_13_port, 
      REGISTERS_21_12_port, REGISTERS_21_11_port, REGISTERS_21_10_port, 
      REGISTERS_21_9_port, REGISTERS_21_8_port, REGISTERS_21_7_port, 
      REGISTERS_21_6_port, REGISTERS_21_5_port, REGISTERS_21_4_port, 
      REGISTERS_21_3_port, REGISTERS_21_2_port, REGISTERS_21_1_port, 
      REGISTERS_21_0_port, REGISTERS_22_63_port, REGISTERS_22_62_port, 
      REGISTERS_22_61_port, REGISTERS_22_60_port, REGISTERS_22_59_port, 
      REGISTERS_22_58_port, REGISTERS_22_57_port, REGISTERS_22_56_port, 
      REGISTERS_22_55_port, REGISTERS_22_54_port, REGISTERS_22_53_port, 
      REGISTERS_22_52_port, REGISTERS_22_51_port, REGISTERS_22_50_port, 
      REGISTERS_22_49_port, REGISTERS_22_48_port, REGISTERS_22_47_port, 
      REGISTERS_22_46_port, REGISTERS_22_45_port, REGISTERS_22_44_port, 
      REGISTERS_22_43_port, REGISTERS_22_42_port, REGISTERS_22_41_port, 
      REGISTERS_22_40_port, REGISTERS_22_39_port, REGISTERS_22_38_port, 
      REGISTERS_22_37_port, REGISTERS_22_36_port, REGISTERS_22_35_port, 
      REGISTERS_22_34_port, REGISTERS_22_33_port, REGISTERS_22_32_port, 
      REGISTERS_22_31_port, REGISTERS_22_30_port, REGISTERS_22_29_port, 
      REGISTERS_22_28_port, REGISTERS_22_27_port, REGISTERS_22_26_port, 
      REGISTERS_22_25_port, REGISTERS_22_24_port, REGISTERS_22_23_port, 
      REGISTERS_22_22_port, REGISTERS_22_21_port, REGISTERS_22_20_port, 
      REGISTERS_22_19_port, REGISTERS_22_18_port, REGISTERS_22_17_port, 
      REGISTERS_22_16_port, REGISTERS_22_15_port, REGISTERS_22_14_port, 
      REGISTERS_22_13_port, REGISTERS_22_12_port, REGISTERS_22_11_port, 
      REGISTERS_22_10_port, REGISTERS_22_9_port, REGISTERS_22_8_port, 
      REGISTERS_22_7_port, REGISTERS_22_6_port, REGISTERS_22_5_port, 
      REGISTERS_22_4_port, REGISTERS_22_3_port, REGISTERS_22_2_port, 
      REGISTERS_22_1_port, REGISTERS_22_0_port, REGISTERS_23_63_port, 
      REGISTERS_23_62_port, REGISTERS_23_61_port, REGISTERS_23_60_port, 
      REGISTERS_23_59_port, REGISTERS_23_58_port, REGISTERS_23_57_port, 
      REGISTERS_23_56_port, REGISTERS_23_55_port, REGISTERS_23_54_port, 
      REGISTERS_23_53_port, REGISTERS_23_52_port, REGISTERS_23_51_port, 
      REGISTERS_23_50_port, REGISTERS_23_49_port, REGISTERS_23_48_port, 
      REGISTERS_23_47_port, REGISTERS_23_46_port, REGISTERS_23_45_port, 
      REGISTERS_23_44_port, REGISTERS_23_43_port, REGISTERS_23_42_port, 
      REGISTERS_23_41_port, REGISTERS_23_40_port, REGISTERS_23_39_port, 
      REGISTERS_23_38_port, REGISTERS_23_37_port, REGISTERS_23_36_port, 
      REGISTERS_23_35_port, REGISTERS_23_34_port, REGISTERS_23_33_port, 
      REGISTERS_23_32_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_63_port, REGISTERS_24_62_port, REGISTERS_24_61_port, 
      REGISTERS_24_60_port, REGISTERS_24_59_port, REGISTERS_24_58_port, 
      REGISTERS_24_57_port, REGISTERS_24_56_port, REGISTERS_24_55_port, 
      REGISTERS_24_54_port, REGISTERS_24_53_port, REGISTERS_24_52_port, 
      REGISTERS_24_51_port, REGISTERS_24_50_port, REGISTERS_24_49_port, 
      REGISTERS_24_48_port, REGISTERS_24_47_port, REGISTERS_24_46_port, 
      REGISTERS_24_45_port, REGISTERS_24_44_port, REGISTERS_24_43_port, 
      REGISTERS_24_42_port, REGISTERS_24_41_port, REGISTERS_24_40_port, 
      REGISTERS_24_39_port, REGISTERS_24_38_port, REGISTERS_24_37_port, 
      REGISTERS_24_36_port, REGISTERS_24_35_port, REGISTERS_24_34_port, 
      REGISTERS_24_33_port, REGISTERS_24_32_port, REGISTERS_24_31_port, 
      REGISTERS_24_30_port, REGISTERS_24_29_port, REGISTERS_24_28_port, 
      REGISTERS_24_27_port, REGISTERS_24_26_port, REGISTERS_24_25_port, 
      REGISTERS_24_24_port, REGISTERS_24_23_port, REGISTERS_24_22_port, 
      REGISTERS_24_21_port, REGISTERS_24_20_port, REGISTERS_24_19_port, 
      REGISTERS_24_18_port, REGISTERS_24_17_port, REGISTERS_24_16_port, 
      REGISTERS_24_15_port, REGISTERS_24_14_port, REGISTERS_24_13_port, 
      REGISTERS_24_12_port, REGISTERS_24_11_port, REGISTERS_24_10_port, 
      REGISTERS_24_9_port, REGISTERS_24_8_port, REGISTERS_24_7_port, 
      REGISTERS_24_6_port, REGISTERS_24_5_port, REGISTERS_24_4_port, 
      REGISTERS_24_3_port, REGISTERS_24_2_port, REGISTERS_24_1_port, 
      REGISTERS_24_0_port, REGISTERS_25_63_port, REGISTERS_25_62_port, 
      REGISTERS_25_61_port, REGISTERS_25_60_port, REGISTERS_25_59_port, 
      REGISTERS_25_58_port, REGISTERS_25_57_port, REGISTERS_25_56_port, 
      REGISTERS_25_55_port, REGISTERS_25_54_port, REGISTERS_25_53_port, 
      REGISTERS_25_52_port, REGISTERS_25_51_port, REGISTERS_25_50_port, 
      REGISTERS_25_49_port, REGISTERS_25_48_port, REGISTERS_25_47_port, 
      REGISTERS_25_46_port, REGISTERS_25_45_port, REGISTERS_25_44_port, 
      REGISTERS_25_43_port, REGISTERS_25_42_port, REGISTERS_25_41_port, 
      REGISTERS_25_40_port, REGISTERS_25_39_port, REGISTERS_25_38_port, 
      REGISTERS_25_37_port, REGISTERS_25_36_port, REGISTERS_25_35_port, 
      REGISTERS_25_34_port, REGISTERS_25_33_port, REGISTERS_25_32_port, 
      REGISTERS_25_31_port, REGISTERS_25_30_port, REGISTERS_25_29_port, 
      REGISTERS_25_28_port, REGISTERS_25_27_port, REGISTERS_25_26_port, 
      REGISTERS_25_25_port, REGISTERS_25_24_port, REGISTERS_25_23_port, 
      REGISTERS_25_22_port, REGISTERS_25_21_port, REGISTERS_25_20_port, 
      REGISTERS_25_19_port, REGISTERS_25_18_port, REGISTERS_25_17_port, 
      REGISTERS_25_16_port, REGISTERS_25_15_port, REGISTERS_25_14_port, 
      REGISTERS_25_13_port, REGISTERS_25_12_port, REGISTERS_25_11_port, 
      REGISTERS_25_10_port, REGISTERS_25_9_port, REGISTERS_25_8_port, 
      REGISTERS_25_7_port, REGISTERS_25_6_port, REGISTERS_25_5_port, 
      REGISTERS_25_4_port, REGISTERS_25_3_port, REGISTERS_25_2_port, 
      REGISTERS_25_1_port, REGISTERS_25_0_port, REGISTERS_26_63_port, 
      REGISTERS_26_62_port, REGISTERS_26_61_port, REGISTERS_26_60_port, 
      REGISTERS_26_59_port, REGISTERS_26_58_port, REGISTERS_26_57_port, 
      REGISTERS_26_56_port, REGISTERS_26_55_port, REGISTERS_26_54_port, 
      REGISTERS_26_53_port, REGISTERS_26_52_port, REGISTERS_26_51_port, 
      REGISTERS_26_50_port, REGISTERS_26_49_port, REGISTERS_26_48_port, 
      REGISTERS_26_47_port, REGISTERS_26_46_port, REGISTERS_26_45_port, 
      REGISTERS_26_44_port, REGISTERS_26_43_port, REGISTERS_26_42_port, 
      REGISTERS_26_41_port, REGISTERS_26_40_port, REGISTERS_26_39_port, 
      REGISTERS_26_38_port, REGISTERS_26_37_port, REGISTERS_26_36_port, 
      REGISTERS_26_35_port, REGISTERS_26_34_port, REGISTERS_26_33_port, 
      REGISTERS_26_32_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_63_port, REGISTERS_27_62_port, REGISTERS_27_61_port, 
      REGISTERS_27_60_port, REGISTERS_27_59_port, REGISTERS_27_58_port, 
      REGISTERS_27_57_port, REGISTERS_27_56_port, REGISTERS_27_55_port, 
      REGISTERS_27_54_port, REGISTERS_27_53_port, REGISTERS_27_52_port, 
      REGISTERS_27_51_port, REGISTERS_27_50_port, REGISTERS_27_49_port, 
      REGISTERS_27_48_port, REGISTERS_27_47_port, REGISTERS_27_46_port, 
      REGISTERS_27_45_port, REGISTERS_27_44_port, REGISTERS_27_43_port, 
      REGISTERS_27_42_port, REGISTERS_27_41_port, REGISTERS_27_40_port, 
      REGISTERS_27_39_port, REGISTERS_27_38_port, REGISTERS_27_37_port, 
      REGISTERS_27_36_port, REGISTERS_27_35_port, REGISTERS_27_34_port, 
      REGISTERS_27_33_port, REGISTERS_27_32_port, REGISTERS_27_31_port, 
      REGISTERS_27_30_port, REGISTERS_27_29_port, REGISTERS_27_28_port, 
      REGISTERS_27_27_port, REGISTERS_27_26_port, REGISTERS_27_25_port, 
      REGISTERS_27_24_port, REGISTERS_27_23_port, REGISTERS_27_22_port, 
      REGISTERS_27_21_port, REGISTERS_27_20_port, REGISTERS_27_19_port, 
      REGISTERS_27_18_port, REGISTERS_27_17_port, REGISTERS_27_16_port, 
      REGISTERS_27_15_port, REGISTERS_27_14_port, REGISTERS_27_13_port, 
      REGISTERS_27_12_port, REGISTERS_27_11_port, REGISTERS_27_10_port, 
      REGISTERS_27_9_port, REGISTERS_27_8_port, REGISTERS_27_7_port, 
      REGISTERS_27_6_port, REGISTERS_27_5_port, REGISTERS_27_4_port, 
      REGISTERS_27_3_port, REGISTERS_27_2_port, REGISTERS_27_1_port, 
      REGISTERS_27_0_port, REGISTERS_28_63_port, REGISTERS_28_62_port, 
      REGISTERS_28_61_port, REGISTERS_28_60_port, REGISTERS_28_59_port, 
      REGISTERS_28_58_port, REGISTERS_28_57_port, REGISTERS_28_56_port, 
      REGISTERS_28_55_port, REGISTERS_28_54_port, REGISTERS_28_53_port, 
      REGISTERS_28_52_port, REGISTERS_28_51_port, REGISTERS_28_50_port, 
      REGISTERS_28_49_port, REGISTERS_28_48_port, REGISTERS_28_47_port, 
      REGISTERS_28_46_port, REGISTERS_28_45_port, REGISTERS_28_44_port, 
      REGISTERS_28_43_port, REGISTERS_28_42_port, REGISTERS_28_41_port, 
      REGISTERS_28_40_port, REGISTERS_28_39_port, REGISTERS_28_38_port, 
      REGISTERS_28_37_port, REGISTERS_28_36_port, REGISTERS_28_35_port, 
      REGISTERS_28_34_port, REGISTERS_28_33_port, REGISTERS_28_32_port, 
      REGISTERS_28_31_port, REGISTERS_28_30_port, REGISTERS_28_29_port, 
      REGISTERS_28_28_port, REGISTERS_28_27_port, REGISTERS_28_26_port, 
      REGISTERS_28_25_port, REGISTERS_28_24_port, REGISTERS_28_23_port, 
      REGISTERS_28_22_port, REGISTERS_28_21_port, REGISTERS_28_20_port, 
      REGISTERS_28_19_port, REGISTERS_28_18_port, REGISTERS_28_17_port, 
      REGISTERS_28_16_port, REGISTERS_28_15_port, REGISTERS_28_14_port, 
      REGISTERS_28_13_port, REGISTERS_28_12_port, REGISTERS_28_11_port, 
      REGISTERS_28_10_port, REGISTERS_28_9_port, REGISTERS_28_8_port, 
      REGISTERS_28_7_port, REGISTERS_28_6_port, REGISTERS_28_5_port, 
      REGISTERS_28_4_port, REGISTERS_28_3_port, REGISTERS_28_2_port, 
      REGISTERS_28_1_port, REGISTERS_28_0_port, REGISTERS_29_63_port, 
      REGISTERS_29_62_port, REGISTERS_29_61_port, REGISTERS_29_60_port, 
      REGISTERS_29_59_port, REGISTERS_29_58_port, REGISTERS_29_57_port, 
      REGISTERS_29_56_port, REGISTERS_29_55_port, REGISTERS_29_54_port, 
      REGISTERS_29_53_port, REGISTERS_29_52_port, REGISTERS_29_51_port, 
      REGISTERS_29_50_port, REGISTERS_29_49_port, REGISTERS_29_48_port, 
      REGISTERS_29_47_port, REGISTERS_29_46_port, REGISTERS_29_45_port, 
      REGISTERS_29_44_port, REGISTERS_29_43_port, REGISTERS_29_42_port, 
      REGISTERS_29_41_port, REGISTERS_29_40_port, REGISTERS_29_39_port, 
      REGISTERS_29_38_port, REGISTERS_29_37_port, REGISTERS_29_36_port, 
      REGISTERS_29_35_port, REGISTERS_29_34_port, REGISTERS_29_33_port, 
      REGISTERS_29_32_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_63_port, REGISTERS_30_62_port, REGISTERS_30_61_port, 
      REGISTERS_30_60_port, REGISTERS_30_59_port, REGISTERS_30_58_port, 
      REGISTERS_30_57_port, REGISTERS_30_56_port, REGISTERS_30_55_port, 
      REGISTERS_30_54_port, REGISTERS_30_53_port, REGISTERS_30_52_port, 
      REGISTERS_30_51_port, REGISTERS_30_50_port, REGISTERS_30_49_port, 
      REGISTERS_30_48_port, REGISTERS_30_47_port, REGISTERS_30_46_port, 
      REGISTERS_30_45_port, REGISTERS_30_44_port, REGISTERS_30_43_port, 
      REGISTERS_30_42_port, REGISTERS_30_41_port, REGISTERS_30_40_port, 
      REGISTERS_30_39_port, REGISTERS_30_38_port, REGISTERS_30_37_port, 
      REGISTERS_30_36_port, REGISTERS_30_35_port, REGISTERS_30_34_port, 
      REGISTERS_30_33_port, REGISTERS_30_32_port, REGISTERS_30_31_port, 
      REGISTERS_30_30_port, REGISTERS_30_29_port, REGISTERS_30_28_port, 
      REGISTERS_30_27_port, REGISTERS_30_26_port, REGISTERS_30_25_port, 
      REGISTERS_30_24_port, REGISTERS_30_23_port, REGISTERS_30_22_port, 
      REGISTERS_30_21_port, REGISTERS_30_20_port, REGISTERS_30_19_port, 
      REGISTERS_30_18_port, REGISTERS_30_17_port, REGISTERS_30_16_port, 
      REGISTERS_30_15_port, REGISTERS_30_14_port, REGISTERS_30_13_port, 
      REGISTERS_30_12_port, REGISTERS_30_11_port, REGISTERS_30_10_port, 
      REGISTERS_30_9_port, REGISTERS_30_8_port, REGISTERS_30_7_port, 
      REGISTERS_30_6_port, REGISTERS_30_5_port, REGISTERS_30_4_port, 
      REGISTERS_30_3_port, REGISTERS_30_2_port, REGISTERS_30_1_port, 
      REGISTERS_30_0_port, REGISTERS_31_63_port, REGISTERS_31_62_port, 
      REGISTERS_31_61_port, REGISTERS_31_60_port, REGISTERS_31_59_port, 
      REGISTERS_31_58_port, REGISTERS_31_57_port, REGISTERS_31_56_port, 
      REGISTERS_31_55_port, REGISTERS_31_54_port, REGISTERS_31_53_port, 
      REGISTERS_31_52_port, REGISTERS_31_51_port, REGISTERS_31_50_port, 
      REGISTERS_31_49_port, REGISTERS_31_48_port, REGISTERS_31_47_port, 
      REGISTERS_31_46_port, REGISTERS_31_45_port, REGISTERS_31_44_port, 
      REGISTERS_31_43_port, REGISTERS_31_42_port, REGISTERS_31_41_port, 
      REGISTERS_31_40_port, REGISTERS_31_39_port, REGISTERS_31_38_port, 
      REGISTERS_31_37_port, REGISTERS_31_36_port, REGISTERS_31_35_port, 
      REGISTERS_31_34_port, REGISTERS_31_33_port, REGISTERS_31_32_port, 
      REGISTERS_31_31_port, REGISTERS_31_30_port, REGISTERS_31_29_port, 
      REGISTERS_31_28_port, REGISTERS_31_27_port, REGISTERS_31_26_port, 
      REGISTERS_31_25_port, REGISTERS_31_24_port, REGISTERS_31_23_port, 
      REGISTERS_31_22_port, REGISTERS_31_21_port, REGISTERS_31_20_port, 
      REGISTERS_31_19_port, REGISTERS_31_18_port, REGISTERS_31_17_port, 
      REGISTERS_31_16_port, REGISTERS_31_15_port, REGISTERS_31_14_port, 
      REGISTERS_31_13_port, REGISTERS_31_12_port, REGISTERS_31_11_port, 
      REGISTERS_31_10_port, REGISTERS_31_9_port, REGISTERS_31_8_port, 
      REGISTERS_31_7_port, REGISTERS_31_6_port, REGISTERS_31_5_port, 
      REGISTERS_31_4_port, REGISTERS_31_3_port, REGISTERS_31_2_port, 
      REGISTERS_31_1_port, REGISTERS_31_0_port, n2456, n2457, n2458, n2459, 
      n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, 
      n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, 
      n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, 
      n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, 
      n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, 
      n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, 
      n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, 
      n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, 
      n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, 
      n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, 
      n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, 
      n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, 
      n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, 
      n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, 
      n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, 
      n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, 
      n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, 
      n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, 
      n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, 
      n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, 
      n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, 
      n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, 
      n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, 
      n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, 
      n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, 
      n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, 
      n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, 
      n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, 
      n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, 
      n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, 
      n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, 
      n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, 
      n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, 
      n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, 
      n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, 
      n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, 
      n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, 
      n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, 
      n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, 
      n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, 
      n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, 
      n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, 
      n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, 
      n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, 
      n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, 
      n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, 
      n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, 
      n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, 
      n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, 
      n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, 
      n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, 
      n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, 
      n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, 
      n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, 
      n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, 
      n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, 
      n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, 
      n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, 
      n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, 
      n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, 
      n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, 
      n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, 
      n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, 
      n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, 
      n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, 
      n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, 
      n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, 
      n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, 
      n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, 
      n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, 
      n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, 
      n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, 
      n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, 
      n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, 
      n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, 
      n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, 
      n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, 
      n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, 
      n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, 
      n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, 
      n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, 
      n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, 
      n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, 
      n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, 
      n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, 
      n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, 
      n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, 
      n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, 
      n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, 
      n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, 
      n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, 
      n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, 
      n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, 
      n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, 
      n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, 
      n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, 
      n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, 
      n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, 
      n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, 
      n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, 
      n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, 
      n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, 
      n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, 
      n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, 
      n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, 
      n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, 
      n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, 
      n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, 
      n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, 
      n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, 
      n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, 
      n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, 
      n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, 
      n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, 
      n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, 
      n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, 
      n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, 
      n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, 
      n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, 
      n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, 
      n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, 
      n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, 
      n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, 
      n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, 
      n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, 
      n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, 
      n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, 
      n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, 
      n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, 
      n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, 
      n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, 
      n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, 
      n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, 
      n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, 
      n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, 
      n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, 
      n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, 
      n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, 
      n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, 
      n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, 
      n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, 
      n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, 
      n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, 
      n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, 
      n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, 
      n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, 
      n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, 
      n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, 
      n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, 
      n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, 
      n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, 
      n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, 
      n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, 
      n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, 
      n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, 
      n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, 
      n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, 
      n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, 
      n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, 
      n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, 
      n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, 
      n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, 
      n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, 
      n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, 
      n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, 
      n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, 
      n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, 
      n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, 
      n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, 
      n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, 
      n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, 
      n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, 
      n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, 
      n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, 
      n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, 
      n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, 
      n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, 
      n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, 
      n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, 
      n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, 
      n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, 
      n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, 
      n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, 
      n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, 
      n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, 
      n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, 
      n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, 
      n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, 
      n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, 
      n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, 
      n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, 
      n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, 
      n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, 
      n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, 
      n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, 
      n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, 
      n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, 
      n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, 
      n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, 
      n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, 
      n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, 
      n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, 
      n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, 
      n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, 
      n4500, n4501, n4502, n4503, n8378, n8379, n8380, n8381, n8382, n8383, 
      n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, 
      n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, 
      n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, 
      n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, 
      n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, 
      n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, 
      n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, 
      n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, 
      n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, 
      n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, 
      n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, 
      n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, 
      n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, 
      n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, 
      n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, 
      n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, 
      n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, 
      n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, 
      n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, 
      n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, 
      n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, 
      n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, 
      n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, 
      n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, 
      n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, 
      n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, 
      n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, 
      n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, 
      n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, 
      n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, 
      n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, 
      n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, 
      n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, 
      n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, 
      n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, 
      n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, 
      n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, 
      n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, 
      n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, 
      n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, 
      n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, 
      n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, 
      n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, 
      n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, 
      n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, 
      n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, 
      n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, 
      n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, 
      n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, 
      n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, 
      n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, 
      n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, 
      n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, 
      n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, 
      n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, 
      n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, 
      n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, 
      n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, 
      n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, 
      n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, 
      n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, 
      n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, 
      n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, 
      n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, 
      n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, 
      n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, 
      n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, 
      n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, 
      n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, 
      n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, 
      n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, 
      n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, 
      n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, 
      n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, 
      n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, 
      n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, 
      n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, 
      n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, 
      n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, 
      n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, 
      n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, 
      n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, 
      n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, 
      n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, 
      n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, 
      n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, 
      n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, 
      n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, 
      n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, 
      n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, 
      n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, 
      n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, 
      n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, 
      n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, 
      n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, 
      n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, 
      n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, 
      n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, 
      n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, 
      n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, 
      n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, 
      n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, 
      n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, 
      n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, 
      n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, 
      n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, 
      n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, 
      n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, 
      n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, 
      n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, 
      n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, 
      n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, 
      n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, 
      n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, 
      n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, 
      n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, 
      n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, 
      n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, 
      n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, 
      n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, 
      n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, 
      n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, 
      n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, 
      n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, 
      n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, 
      n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, 
      n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, 
      n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, 
      n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, 
      n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, 
      n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, 
      n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, 
      n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, 
      n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, 
      n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, 
      n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, 
      n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, 
      n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, 
      n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, 
      n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, 
      n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, 
      n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, 
      n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, 
      n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, 
      n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, 
      n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, 
      n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, 
      n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, 
      n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, 
      n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, 
      n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, 
      n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, 
      n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, 
      n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, 
      n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, 
      n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, 
      n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, 
      n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, 
      n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, 
      n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, 
      n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, 
      n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, 
      n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, 
      n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, 
      n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, 
      n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, 
      n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, 
      n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, 
      n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, 
      n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, 
      n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, 
      n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, 
      n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, 
      n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, 
      n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, 
      n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, 
      n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, 
      n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, 
      n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, 
      n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, 
      n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, 
      n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, 
      n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, 
      n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, 
      n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, 
      n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, 
      n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, 
      n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, 
      n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, 
      n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, 
      n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, 
      n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, 
      n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, 
      n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, 
      n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, 
      n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, 
      n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, 
      n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, 
      n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, 
      n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, 
      n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, 
      n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, 
      n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, 
      n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, 
      n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, 
      n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, 
      n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, 
      n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, 
      n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, 
      n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, 
      n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, 
      n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, 
      n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, 
      n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, 
      n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, 
      n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, 
      n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, 
      n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, 
      n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, 
      n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, 
      n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, 
      n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, 
      n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, 
      n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, 
      n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, 
      n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, 
      n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, 
      n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, 
      n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, 
      n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, 
      n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, 
      n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, 
      n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, 
      n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, 
      n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, 
      n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, 
      n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, 
      n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, 
      n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, 
      n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, 
      n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, 
      n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, 
      n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, 
      n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, 
      n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, 
      n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, 
      n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, 
      n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, 
      n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, 
      n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, 
      n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, 
      n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, 
      n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, 
      n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, 
      n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, 
      n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, 
      n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, 
      n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, 
      n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, 
      n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, 
      n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, 
      n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, 
      n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, 
      n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, 
      n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, 
      n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, 
      n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, 
      n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, 
      n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, 
      n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, 
      n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, 
      n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, 
      n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, 
      n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, 
      n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, 
      n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, 
      n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, 
      n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, 
      n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, 
      n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, 
      n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, 
      n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, 
      n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, 
      n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, 
      n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, 
      n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, 
      n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, 
      n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, 
      n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, 
      n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, 
      n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, 
      n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, 
      n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, 
      n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, 
      n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, 
      n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, 
      n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, 
      n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, 
      n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, 
      n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, 
      n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, 
      n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, 
      n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, 
      n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, 
      n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, 
      n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, 
      n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, 
      n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, 
      n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, 
      n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, 
      n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, 
      n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, 
      n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, 
      n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, 
      n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, 
      n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, 
      n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, 
      n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, 
      n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, 
      n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, 
      n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, 
      n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, 
      n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, 
      n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, 
      n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, 
      n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, 
      n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, 
      n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, 
      n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, 
      n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, 
      n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, 
      n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, 
      n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, 
      n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, 
      n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, 
      n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, 
      n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, 
      n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, 
      n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, 
      n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, 
      n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, 
      n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, 
      n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, 
      n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, 
      n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, 
      n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, 
      n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, 
      n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, 
      n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, 
      n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, 
      n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, 
      n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, 
      n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, 
      n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, 
      n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, 
      n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, 
      n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, 
      n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, 
      n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, 
      n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, 
      n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, 
      n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, 
      n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, 
      n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, 
      n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, 
      n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, 
      n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, 
      n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, 
      n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, 
      n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, 
      n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, 
      n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, 
      n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, 
      n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, 
      n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, 
      n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, 
      n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, 
      n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, 
      n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, 
      n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, 
      n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, 
      n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, 
      n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, 
      n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, 
      n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, 
      n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, 
      n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, 
      n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, 
      n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, 
      n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, 
      n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, 
      n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, 
      n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, 
      n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, 
      n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, 
      n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, 
      n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, 
      n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, 
      n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, 
      n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, 
      n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, 
      n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, 
      n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, 
      n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, 
      n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, 
      n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, 
      n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, 
      n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, 
      n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, 
      n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, 
      n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, 
      n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, 
      n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, 
      n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, 
      n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, 
      n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, 
      n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, 
      n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, 
      n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, 
      n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, 
      n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, 
      n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, 
      n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, 
      n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, 
      n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, 
      n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, 
      n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, 
      n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, 
      n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, 
      n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, 
      n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, 
      n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, 
      n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, 
      n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, 
      n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, 
      n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, 
      n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, 
      n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, 
      n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, 
      n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, 
      n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, 
      n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, 
      n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, 
      n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, 
      n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, 
      n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, 
      n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, 
      n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, 
      n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, 
      n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, 
      n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, 
      n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, 
      n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, 
      n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, 
      n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, 
      n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, 
      n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, 
      n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, 
      n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, 
      n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, 
      n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, 
      n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, 
      n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, 
      n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, 
      n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, 
      n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, 
      n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, 
      n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, 
      n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, 
      n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, 
      n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, 
      n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, 
      n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, 
      n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, 
      n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, 
      n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, 
      n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, 
      n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, 
      n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, 
      n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, 
      n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, 
      n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, 
      n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, 
      n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, 
      n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, 
      n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, 
      n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, 
      n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, 
      n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, 
      n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, 
      n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, 
      n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, 
      n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, 
      n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, 
      n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, 
      n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, 
      n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, 
      n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, 
      n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, 
      n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, 
      n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, 
      n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, 
      n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, 
      n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, 
      n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, 
      n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, 
      n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, 
      n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, 
      n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, 
      n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, 
      n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, 
      n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, 
      n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, 
      n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, 
      n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, 
      n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, 
      n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, 
      n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, 
      n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, 
      n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, 
      n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, 
      n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, 
      n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, 
      n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, 
      n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, 
      n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, 
      n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, 
      n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, 
      n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, 
      n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, 
      n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, 
      n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, 
      n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, 
      n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, 
      n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, 
      n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, 
      n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, 
      n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, 
      n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, 
      n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, 
      n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, 
      n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, 
      n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, 
      n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, 
      n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, 
      n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, 
      n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, 
      n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, 
      n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, 
      n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, 
      n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, 
      n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, 
      n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, 
      n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, 
      n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, 
      n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, 
      n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, 
      n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, 
      n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, 
      n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, 
      n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, 
      n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, 
      n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, 
      n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, 
      n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, 
      n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, 
      n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, 
      n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, 
      n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, 
      n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, 
      n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, 
      n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, 
      n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, 
      n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, 
      n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, 
      n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, 
      n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, 
      n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, 
      n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, 
      n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, 
      n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, 
      n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, 
      n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, 
      n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, 
      n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, 
      n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, 
      n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, 
      n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, 
      n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, 
      n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, 
      n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, 
      n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, 
      n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, 
      n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, 
      n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, 
      n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, 
      n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, 
      n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, 
      n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, 
      n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, 
      n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, 
      n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, 
      n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930 : 
      std_logic;

begin
   
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n4503, CK => CLK, Q => 
                           REGISTERS_0_63_port, QN => n16884);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n4502, CK => CLK, Q => 
                           REGISTERS_0_62_port, QN => n18017);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n4501, CK => CLK, Q => 
                           REGISTERS_0_61_port, QN => n18243);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n4500, CK => CLK, Q => 
                           REGISTERS_0_60_port, QN => n18018);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n4499, CK => CLK, Q => 
                           REGISTERS_0_59_port, QN => n18244);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n4498, CK => CLK, Q => 
                           REGISTERS_0_58_port, QN => n18019);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n4497, CK => CLK, Q => 
                           REGISTERS_0_57_port, QN => n18020);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n4496, CK => CLK, Q => 
                           REGISTERS_0_56_port, QN => n18245);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n4495, CK => CLK, Q => 
                           REGISTERS_0_55_port, QN => n18246);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n4494, CK => CLK, Q => 
                           REGISTERS_0_54_port, QN => n18021);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n4493, CK => CLK, Q => 
                           REGISTERS_0_53_port, QN => n18247);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n4492, CK => CLK, Q => 
                           REGISTERS_0_52_port, QN => n18248);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n4491, CK => CLK, Q => 
                           REGISTERS_0_51_port, QN => n18022);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n4490, CK => CLK, Q => 
                           REGISTERS_0_50_port, QN => n18023);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n4489, CK => CLK, Q => 
                           REGISTERS_0_49_port, QN => n18024);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n4488, CK => CLK, Q => 
                           REGISTERS_0_48_port, QN => n18249);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n4487, CK => CLK, Q => 
                           REGISTERS_0_47_port, QN => n17388);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n4486, CK => CLK, Q => 
                           REGISTERS_0_46_port, QN => n17172);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n4485, CK => CLK, Q => 
                           REGISTERS_0_45_port, QN => n17389);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n4484, CK => CLK, Q => 
                           REGISTERS_0_44_port, QN => n17173);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n4483, CK => CLK, Q => 
                           REGISTERS_0_43_port, QN => n17390);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n4482, CK => CLK, Q => 
                           REGISTERS_0_42_port, QN => n17174);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n4481, CK => CLK, Q => 
                           REGISTERS_0_41_port, QN => n17175);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n4480, CK => CLK, Q => 
                           REGISTERS_0_40_port, QN => n17176);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n4479, CK => CLK, Q => 
                           REGISTERS_0_39_port, QN => n17177);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n4478, CK => CLK, Q => 
                           REGISTERS_0_38_port, QN => n17178);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n4477, CK => CLK, Q => 
                           REGISTERS_0_37_port, QN => n17179);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n4476, CK => CLK, Q => 
                           REGISTERS_0_36_port, QN => n17391);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n4475, CK => CLK, Q => 
                           REGISTERS_0_35_port, QN => n18025);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n4474, CK => CLK, Q => 
                           REGISTERS_0_34_port, QN => n18250);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n4473, CK => CLK, Q => 
                           REGISTERS_0_33_port, QN => n18026);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n4472, CK => CLK, Q => 
                           REGISTERS_0_32_port, QN => n18027);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n4471, CK => CLK, Q => 
                           REGISTERS_0_31_port, QN => n18251);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n4470, CK => CLK, Q => 
                           REGISTERS_0_30_port, QN => n18252);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n4469, CK => CLK, Q => 
                           REGISTERS_0_29_port, QN => n18253);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n4468, CK => CLK, Q => 
                           REGISTERS_0_28_port, QN => n18254);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n4467, CK => CLK, Q => 
                           REGISTERS_0_27_port, QN => n17180);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n4466, CK => CLK, Q => 
                           REGISTERS_0_26_port, QN => n17392);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n4465, CK => CLK, Q => 
                           REGISTERS_0_25_port, QN => n17393);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n4464, CK => CLK, Q => 
                           REGISTERS_0_24_port, QN => n17394);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n4463, CK => CLK, Q => 
                           REGISTERS_0_23_port, QN => n17181);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n4462, CK => CLK, Q => 
                           REGISTERS_0_22_port, QN => n17182);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n4461, CK => CLK, Q => 
                           REGISTERS_0_21_port, QN => n17395);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n4460, CK => CLK, Q => 
                           REGISTERS_0_20_port, QN => n17183);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n4459, CK => CLK, Q => 
                           REGISTERS_0_19_port, QN => n17184);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n4458, CK => CLK, Q => 
                           REGISTERS_0_18_port, QN => n17396);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n4457, CK => CLK, Q => 
                           REGISTERS_0_17_port, QN => n17185);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n4456, CK => CLK, Q => 
                           REGISTERS_0_16_port, QN => n17397);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n4455, CK => CLK, Q => 
                           REGISTERS_0_15_port, QN => n18028);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n4454, CK => CLK, Q => 
                           REGISTERS_0_14_port, QN => n18029);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n4453, CK => CLK, Q => 
                           REGISTERS_0_13_port, QN => n18255);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n4452, CK => CLK, Q => 
                           REGISTERS_0_12_port, QN => n17398);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n4451, CK => CLK, Q => 
                           REGISTERS_0_11_port, QN => n17399);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n4450, CK => CLK, Q => 
                           REGISTERS_0_10_port, QN => n17186);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n4449, CK => CLK, Q => 
                           REGISTERS_0_9_port, QN => n17187);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n4448, CK => CLK, Q => 
                           REGISTERS_0_8_port, QN => n17188);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n4447, CK => CLK, Q => 
                           REGISTERS_0_7_port, QN => n17400);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n4446, CK => CLK, Q => 
                           REGISTERS_0_6_port, QN => n17189);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n4445, CK => CLK, Q => 
                           REGISTERS_0_5_port, QN => n17401);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n4444, CK => CLK, Q => 
                           REGISTERS_0_4_port, QN => n17402);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n4443, CK => CLK, Q => 
                           REGISTERS_0_3_port, QN => n17403);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n4442, CK => CLK, Q => 
                           REGISTERS_0_2_port, QN => n17404);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n4441, CK => CLK, Q => 
                           REGISTERS_0_1_port, QN => n17405);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n4440, CK => CLK, Q => 
                           REGISTERS_0_0_port, QN => n18256);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n4439, CK => CLK, Q => 
                           REGISTERS_1_63_port, QN => n17105);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n4438, CK => CLK, Q => 
                           REGISTERS_1_62_port, QN => n18257);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n4437, CK => CLK, Q => 
                           REGISTERS_1_61_port, QN => n18701);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n4436, CK => CLK, Q => 
                           REGISTERS_1_60_port, QN => n18258);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n4435, CK => CLK, Q => 
                           REGISTERS_1_59_port, QN => n18702);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n4434, CK => CLK, Q => 
                           REGISTERS_1_58_port, QN => n18259);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n4433, CK => CLK, Q => 
                           REGISTERS_1_57_port, QN => n18703);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n4432, CK => CLK, Q => 
                           REGISTERS_1_56_port, QN => n18260);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n4431, CK => CLK, Q => 
                           REGISTERS_1_55_port, QN => n18030);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n4430, CK => CLK, Q => 
                           REGISTERS_1_54_port, QN => n18704);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n4429, CK => CLK, Q => 
                           REGISTERS_1_53_port, QN => n18261);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n4428, CK => CLK, Q => 
                           REGISTERS_1_52_port, QN => n18262);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n4427, CK => CLK, Q => 
                           REGISTERS_1_51_port, QN => n18263);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n4426, CK => CLK, Q => 
                           REGISTERS_1_50_port, QN => n18705);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n4425, CK => CLK, Q => 
                           REGISTERS_1_49_port, QN => n18706);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n4424, CK => CLK, Q => 
                           REGISTERS_1_48_port, QN => n18707);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n4423, CK => CLK, Q => 
                           REGISTERS_1_47_port, QN => n18264);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n4422, CK => CLK, Q => 
                           REGISTERS_1_46_port, QN => n18265);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n4421, CK => CLK, Q => 
                           REGISTERS_1_45_port, QN => n18708);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n4420, CK => CLK, Q => 
                           REGISTERS_1_44_port, QN => n18266);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n4419, CK => CLK, Q => 
                           REGISTERS_1_43_port, QN => n18267);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n4418, CK => CLK, Q => 
                           REGISTERS_1_42_port, QN => n18709);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n4417, CK => CLK, Q => 
                           REGISTERS_1_41_port, QN => n18268);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n4416, CK => CLK, Q => 
                           REGISTERS_1_40_port, QN => n18031);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n4415, CK => CLK, Q => 
                           REGISTERS_1_39_port, QN => n18269);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n4414, CK => CLK, Q => 
                           REGISTERS_1_38_port, QN => n18270);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n4413, CK => CLK, Q => 
                           REGISTERS_1_37_port, QN => n18271);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n4412, CK => CLK, Q => 
                           REGISTERS_1_36_port, QN => n18272);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n4411, CK => CLK, Q => 
                           REGISTERS_1_35_port, QN => n18710);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n4410, CK => CLK, Q => 
                           REGISTERS_1_34_port, QN => n18273);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n4409, CK => CLK, Q => 
                           REGISTERS_1_33_port, QN => n18274);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n4408, CK => CLK, Q => 
                           REGISTERS_1_32_port, QN => n18275);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n4407, CK => CLK, Q => 
                           REGISTERS_1_31_port, QN => n18032);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n4406, CK => CLK, Q => 
                           REGISTERS_1_30_port, QN => n18711);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n4405, CK => CLK, Q => 
                           REGISTERS_1_29_port, QN => n18276);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n4404, CK => n13730, Q => 
                           REGISTERS_1_28_port, QN => n18277);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n4403, CK => CLK, Q => 
                           REGISTERS_1_27_port, QN => n17794);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n4402, CK => CLK, Q => 
                           REGISTERS_1_26_port, QN => n17406);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n4401, CK => CLK, Q => 
                           REGISTERS_1_25_port, QN => n17795);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n4400, CK => CLK, Q => 
                           REGISTERS_1_24_port, QN => n17407);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n4399, CK => CLK, Q => 
                           REGISTERS_1_23_port, QN => n17796);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n4398, CK => CLK, Q => 
                           REGISTERS_1_22_port, QN => n17408);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n4397, CK => CLK, Q => 
                           REGISTERS_1_21_port, QN => n17190);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n4396, CK => CLK, Q => 
                           REGISTERS_1_20_port, QN => n17191);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n4395, CK => CLK, Q => 
                           REGISTERS_1_19_port, QN => n17409);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n4394, CK => CLK, Q => 
                           REGISTERS_1_18_port, QN => n17797);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n4393, CK => CLK, Q => 
                           REGISTERS_1_17_port, QN => n17798);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n4392, CK => CLK, Q => 
                           REGISTERS_1_16_port, QN => n17799);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n4391, CK => CLK, Q => 
                           REGISTERS_1_15_port, QN => n18712);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n4390, CK => CLK, Q => 
                           REGISTERS_1_14_port, QN => n18713);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n4389, CK => CLK, Q => 
                           REGISTERS_1_13_port, QN => n18714);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n4388, CK => CLK, Q => 
                           REGISTERS_1_12_port, QN => n18278);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n4387, CK => CLK, Q => 
                           REGISTERS_1_11_port, QN => n18715);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n4386, CK => CLK, Q => 
                           REGISTERS_1_10_port, QN => n18033);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n4385, CK => CLK, Q => 
                           REGISTERS_1_9_port, QN => n18279);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n4384, CK => CLK, Q => 
                           REGISTERS_1_8_port, QN => n18280);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n4383, CK => CLK, Q => 
                           REGISTERS_1_7_port, QN => n18281);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n4382, CK => CLK, Q => 
                           REGISTERS_1_6_port, QN => n18282);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n4381, CK => CLK, Q => 
                           REGISTERS_1_5_port, QN => n18283);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n4380, CK => CLK, Q => 
                           REGISTERS_1_4_port, QN => n18716);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n4379, CK => CLK, Q => 
                           REGISTERS_1_3_port, QN => n18717);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n4378, CK => CLK, Q => 
                           REGISTERS_1_2_port, QN => n18284);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n4377, CK => CLK, Q => 
                           REGISTERS_1_1_port, QN => n18718);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n4376, CK => CLK, Q => 
                           REGISTERS_1_0_port, QN => n18719);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n4375, CK => CLK, Q => 
                           REGISTERS_2_63_port, QN => n17106);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n4374, CK => CLK, Q => 
                           REGISTERS_2_62_port, QN => n18720);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n4373, CK => CLK, Q => 
                           REGISTERS_2_61_port, QN => n18285);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n4372, CK => CLK, Q => 
                           REGISTERS_2_60_port, QN => n18721);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n4371, CK => CLK, Q => 
                           REGISTERS_2_59_port, QN => n18722);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n4370, CK => CLK, Q => 
                           REGISTERS_2_58_port, QN => n18723);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n4369, CK => CLK, Q => 
                           REGISTERS_2_57_port, QN => n18286);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n4368, CK => CLK, Q => 
                           REGISTERS_2_56_port, QN => n18287);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n4367, CK => CLK, Q => 
                           REGISTERS_2_55_port, QN => n18288);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n4366, CK => CLK, Q => 
                           REGISTERS_2_54_port, QN => n18724);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n4365, CK => CLK, Q => 
                           REGISTERS_2_53_port, QN => n18725);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n4364, CK => CLK, Q => 
                           REGISTERS_2_52_port, QN => n18289);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n4363, CK => CLK, Q => 
                           REGISTERS_2_51_port, QN => n18726);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n4362, CK => CLK, Q => 
                           REGISTERS_2_50_port, QN => n18727);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n4361, CK => CLK, Q => 
                           REGISTERS_2_49_port, QN => n18290);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n4360, CK => CLK, Q => 
                           REGISTERS_2_48_port, QN => n18728);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n4359, CK => CLK, Q => 
                           REGISTERS_2_47_port, QN => n18291);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n4358, CK => n13730, Q => 
                           REGISTERS_2_46_port, QN => n18729);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n4357, CK => CLK, Q => 
                           REGISTERS_2_45_port, QN => n18730);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n4356, CK => CLK, Q => 
                           REGISTERS_2_44_port, QN => n18731);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n4355, CK => CLK, Q => 
                           REGISTERS_2_43_port, QN => n18732);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n4354, CK => CLK, Q => 
                           REGISTERS_2_42_port, QN => n18292);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n4353, CK => CLK, Q => 
                           REGISTERS_2_41_port, QN => n18293);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n4352, CK => CLK, Q => 
                           REGISTERS_2_40_port, QN => n18733);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n4351, CK => CLK, Q => 
                           REGISTERS_2_39_port, QN => n18734);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n4350, CK => CLK, Q => 
                           REGISTERS_2_38_port, QN => n18735);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n4349, CK => CLK, Q => 
                           REGISTERS_2_37_port, QN => n18736);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n4348, CK => CLK, Q => 
                           REGISTERS_2_36_port, QN => n18294);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n4347, CK => CLK, Q => 
                           REGISTERS_2_35_port, QN => n18295);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n4346, CK => CLK, Q => 
                           REGISTERS_2_34_port, QN => n18737);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n4345, CK => CLK, Q => 
                           REGISTERS_2_33_port, QN => n18738);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n4344, CK => CLK, Q => 
                           REGISTERS_2_32_port, QN => n18296);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n4343, CK => CLK, Q => 
                           REGISTERS_2_31_port, QN => n18297);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n4342, CK => CLK, Q => 
                           REGISTERS_2_30_port, QN => n18298);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n4341, CK => CLK, Q => 
                           REGISTERS_2_29_port, QN => n18299);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n4340, CK => CLK, Q => 
                           REGISTERS_2_28_port, QN => n18300);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n4339, CK => CLK, Q => 
                           REGISTERS_2_27_port, QN => n17800);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n4338, CK => CLK, Q => 
                           REGISTERS_2_26_port, QN => n17801);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n4337, CK => CLK, Q => 
                           REGISTERS_2_25_port, QN => n17410);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n4336, CK => CLK, Q => 
                           REGISTERS_2_24_port, QN => n17411);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n4335, CK => CLK, Q => 
                           REGISTERS_2_23_port, QN => n17412);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n4334, CK => CLK, Q => 
                           REGISTERS_2_22_port, QN => n17802);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n4333, CK => CLK, Q => 
                           REGISTERS_2_21_port, QN => n17803);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n4332, CK => CLK, Q => 
                           REGISTERS_2_20_port, QN => n17804);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n4331, CK => CLK, Q => 
                           REGISTERS_2_19_port, QN => n17805);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n4330, CK => CLK, Q => 
                           REGISTERS_2_18_port, QN => n17806);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n4329, CK => CLK, Q => 
                           REGISTERS_2_17_port, QN => n17413);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n4328, CK => CLK, Q => 
                           REGISTERS_2_16_port, QN => n17414);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n4327, CK => CLK, Q => 
                           REGISTERS_2_15_port, QN => n18301);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n4326, CK => CLK, Q => 
                           REGISTERS_2_14_port, QN => n18739);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n4325, CK => CLK, Q => 
                           REGISTERS_2_13_port, QN => n18302);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n4324, CK => CLK, Q => 
                           REGISTERS_2_12_port, QN => n18303);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n4323, CK => CLK, Q => 
                           REGISTERS_2_11_port, QN => n18740);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n4322, CK => CLK, Q => 
                           REGISTERS_2_10_port, QN => n18304);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n4321, CK => CLK, Q => 
                           REGISTERS_2_9_port, QN => n18741);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n4320, CK => CLK, Q => 
                           REGISTERS_2_8_port, QN => n18742);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n4319, CK => CLK, Q => 
                           REGISTERS_2_7_port, QN => n18305);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n4318, CK => CLK, Q => 
                           REGISTERS_2_6_port, QN => n18743);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n4317, CK => CLK, Q => 
                           REGISTERS_2_5_port, QN => n18306);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n4316, CK => CLK, Q => 
                           REGISTERS_2_4_port, QN => n18744);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n4315, CK => CLK, Q => 
                           REGISTERS_2_3_port, QN => n18307);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n4314, CK => CLK, Q => 
                           REGISTERS_2_2_port, QN => n18308);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n4313, CK => CLK, Q => 
                           REGISTERS_2_1_port, QN => n18309);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n4312, CK => CLK, Q => 
                           REGISTERS_2_0_port, QN => n18310);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n4311, CK => CLK, Q => 
                           REGISTERS_3_63_port, QN => n16963);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n4310, CK => CLK, Q => 
                           REGISTERS_3_62_port, QN => n18311);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n4309, CK => CLK, Q => 
                           REGISTERS_3_61_port, QN => n18034);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n4308, CK => CLK, Q => 
                           REGISTERS_3_60_port, QN => n18312);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n4307, CK => CLK, Q => 
                           REGISTERS_3_59_port, QN => n18313);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n4306, CK => CLK, Q => 
                           REGISTERS_3_58_port, QN => n18314);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n4305, CK => CLK, Q => 
                           REGISTERS_3_57_port, QN => n18315);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n4304, CK => CLK, Q => 
                           REGISTERS_3_56_port, QN => n18035);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n4303, CK => CLK, Q => 
                           REGISTERS_3_55_port, QN => n18745);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n4302, CK => CLK, Q => 
                           REGISTERS_3_54_port, QN => n18316);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n4301, CK => CLK, Q => 
                           REGISTERS_3_53_port, QN => n18317);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n4300, CK => CLK, Q => 
                           REGISTERS_3_52_port, QN => n18746);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n4299, CK => CLK, Q => 
                           REGISTERS_3_51_port, QN => n18747);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n4298, CK => CLK, Q => 
                           REGISTERS_3_50_port, QN => n18318);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n4297, CK => CLK, Q => 
                           REGISTERS_3_49_port, QN => n18319);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n4296, CK => CLK, Q => 
                           REGISTERS_3_48_port, QN => n18036);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n4295, CK => CLK, Q => 
                           REGISTERS_3_47_port, QN => n18320);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n4294, CK => CLK, Q => 
                           REGISTERS_3_46_port, QN => n18321);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n4293, CK => CLK, Q => 
                           REGISTERS_3_45_port, QN => n18322);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n4292, CK => CLK, Q => 
                           REGISTERS_3_44_port, QN => n18323);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n4291, CK => CLK, Q => 
                           REGISTERS_3_43_port, QN => n18324);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n4290, CK => CLK, Q => 
                           REGISTERS_3_42_port, QN => n18325);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n4289, CK => CLK, Q => 
                           REGISTERS_3_41_port, QN => n18326);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n4288, CK => CLK, Q => 
                           REGISTERS_3_40_port, QN => n18327);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n4287, CK => CLK, Q => 
                           REGISTERS_3_39_port, QN => n18328);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n4286, CK => CLK, Q => 
                           REGISTERS_3_38_port, QN => n18748);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n4285, CK => CLK, Q => 
                           REGISTERS_3_37_port, QN => n18329);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n4284, CK => CLK, Q => 
                           REGISTERS_3_36_port, QN => n18749);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n4283, CK => CLK, Q => 
                           REGISTERS_3_35_port, QN => n18750);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n4282, CK => CLK, Q => 
                           REGISTERS_3_34_port, QN => n18330);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n4281, CK => CLK, Q => 
                           REGISTERS_3_33_port, QN => n18037);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n4280, CK => CLK, Q => 
                           REGISTERS_3_32_port, QN => n18751);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n4279, CK => CLK, Q => 
                           REGISTERS_3_31_port, QN => n18331);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n4278, CK => CLK, Q => 
                           REGISTERS_3_30_port, QN => n18332);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n4277, CK => CLK, Q => 
                           REGISTERS_3_29_port, QN => n18752);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n4276, CK => CLK, Q => 
                           REGISTERS_3_28_port, QN => n18753);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n4275, CK => CLK, Q => 
                           REGISTERS_3_27_port, QN => n17415);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n4274, CK => CLK, Q => 
                           REGISTERS_3_26_port, QN => n17416);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n4273, CK => CLK, Q => 
                           REGISTERS_3_25_port, QN => n17192);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n4272, CK => CLK, Q => 
                           REGISTERS_3_24_port, QN => n17807);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n4271, CK => CLK, Q => 
                           REGISTERS_3_23_port, QN => n17808);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n4270, CK => CLK, Q => 
                           REGISTERS_3_22_port, QN => n17417);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n4269, CK => CLK, Q => 
                           REGISTERS_3_21_port, QN => n17418);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n4268, CK => CLK, Q => 
                           REGISTERS_3_20_port, QN => n17193);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n4267, CK => CLK, Q => 
                           REGISTERS_3_19_port, QN => n17419);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n4266, CK => CLK, Q => 
                           REGISTERS_3_18_port, QN => n17420);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n4265, CK => CLK, Q => 
                           REGISTERS_3_17_port, QN => n17809);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n4264, CK => CLK, Q => 
                           REGISTERS_3_16_port, QN => n17421);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n4263, CK => CLK, Q => 
                           REGISTERS_3_15_port, QN => n18754);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n4262, CK => CLK, Q => 
                           REGISTERS_3_14_port, QN => n18038);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n4261, CK => CLK, Q => 
                           REGISTERS_3_13_port, QN => n18039);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n4260, CK => CLK, Q => 
                           REGISTERS_3_12_port, QN => n18755);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n4259, CK => CLK, Q => 
                           REGISTERS_3_11_port, QN => n18333);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n4258, CK => CLK, Q => 
                           REGISTERS_3_10_port, QN => n18334);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n4257, CK => CLK, Q => 
                           REGISTERS_3_9_port, QN => n18040);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n4256, CK => CLK, Q => 
                           REGISTERS_3_8_port, QN => n18335);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n4255, CK => CLK, Q => 
                           REGISTERS_3_7_port, QN => n18041);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n4254, CK => CLK, Q => 
                           REGISTERS_3_6_port, QN => n18042);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n4253, CK => CLK, Q => 
                           REGISTERS_3_5_port, QN => n18756);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n4252, CK => CLK, Q => 
                           REGISTERS_3_4_port, QN => n18336);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n4251, CK => CLK, Q => 
                           REGISTERS_3_3_port, QN => n18337);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n4250, CK => CLK, Q => 
                           REGISTERS_3_2_port, QN => n18757);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n4249, CK => CLK, Q => 
                           REGISTERS_3_1_port, QN => n18043);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n4248, CK => CLK, Q => 
                           REGISTERS_3_0_port, QN => n18044);
   REGISTERS_reg_4_63_inst : DFF_X1 port map( D => n4247, CK => n13730, Q => 
                           REGISTERS_4_63_port, QN => n16885);
   REGISTERS_reg_4_62_inst : DFF_X1 port map( D => n4246, CK => CLK, Q => 
                           REGISTERS_4_62_port, QN => n18338);
   REGISTERS_reg_4_61_inst : DFF_X1 port map( D => n4245, CK => CLK, Q => 
                           REGISTERS_4_61_port, QN => n18045);
   REGISTERS_reg_4_60_inst : DFF_X1 port map( D => n4244, CK => CLK, Q => 
                           REGISTERS_4_60_port, QN => n18339);
   REGISTERS_reg_4_59_inst : DFF_X1 port map( D => n4243, CK => CLK, Q => 
                           REGISTERS_4_59_port, QN => n18046);
   REGISTERS_reg_4_58_inst : DFF_X1 port map( D => n4242, CK => CLK, Q => 
                           REGISTERS_4_58_port, QN => n18340);
   REGISTERS_reg_4_57_inst : DFF_X1 port map( D => n4241, CK => CLK, Q => 
                           REGISTERS_4_57_port, QN => n18341);
   REGISTERS_reg_4_56_inst : DFF_X1 port map( D => n4240, CK => CLK, Q => 
                           REGISTERS_4_56_port, QN => n18047);
   REGISTERS_reg_4_55_inst : DFF_X1 port map( D => n4239, CK => CLK, Q => 
                           REGISTERS_4_55_port, QN => n18048);
   REGISTERS_reg_4_54_inst : DFF_X1 port map( D => n4238, CK => CLK, Q => 
                           REGISTERS_4_54_port, QN => n18342);
   REGISTERS_reg_4_53_inst : DFF_X1 port map( D => n4237, CK => CLK, Q => 
                           REGISTERS_4_53_port, QN => n18343);
   REGISTERS_reg_4_52_inst : DFF_X1 port map( D => n4236, CK => CLK, Q => 
                           REGISTERS_4_52_port, QN => n18049);
   REGISTERS_reg_4_51_inst : DFF_X1 port map( D => n4235, CK => CLK, Q => 
                           REGISTERS_4_51_port, QN => n18050);
   REGISTERS_reg_4_50_inst : DFF_X1 port map( D => n4234, CK => CLK, Q => 
                           REGISTERS_4_50_port, QN => n18051);
   REGISTERS_reg_4_49_inst : DFF_X1 port map( D => n4233, CK => CLK, Q => 
                           REGISTERS_4_49_port, QN => n18052);
   REGISTERS_reg_4_48_inst : DFF_X1 port map( D => n4232, CK => CLK, Q => 
                           REGISTERS_4_48_port, QN => n18053);
   REGISTERS_reg_4_47_inst : DFF_X1 port map( D => n4231, CK => CLK, Q => 
                           REGISTERS_4_47_port, QN => n18758);
   REGISTERS_reg_4_46_inst : DFF_X1 port map( D => n4230, CK => CLK, Q => 
                           REGISTERS_4_46_port, QN => n18054);
   REGISTERS_reg_4_45_inst : DFF_X1 port map( D => n4229, CK => CLK, Q => 
                           REGISTERS_4_45_port, QN => n18055);
   REGISTERS_reg_4_44_inst : DFF_X1 port map( D => n4228, CK => CLK, Q => 
                           REGISTERS_4_44_port, QN => n18344);
   REGISTERS_reg_4_43_inst : DFF_X1 port map( D => n4227, CK => CLK, Q => 
                           REGISTERS_4_43_port, QN => n18056);
   REGISTERS_reg_4_42_inst : DFF_X1 port map( D => n4226, CK => CLK, Q => 
                           REGISTERS_4_42_port, QN => n18057);
   REGISTERS_reg_4_41_inst : DFF_X1 port map( D => n4225, CK => CLK, Q => 
                           REGISTERS_4_41_port, QN => n18345);
   REGISTERS_reg_4_40_inst : DFF_X1 port map( D => n4224, CK => CLK, Q => 
                           REGISTERS_4_40_port, QN => n18058);
   REGISTERS_reg_4_39_inst : DFF_X1 port map( D => n4223, CK => CLK, Q => 
                           REGISTERS_4_39_port, QN => n18346);
   REGISTERS_reg_4_38_inst : DFF_X1 port map( D => n4222, CK => CLK, Q => 
                           REGISTERS_4_38_port, QN => n18347);
   REGISTERS_reg_4_37_inst : DFF_X1 port map( D => n4221, CK => CLK, Q => 
                           REGISTERS_4_37_port, QN => n18348);
   REGISTERS_reg_4_36_inst : DFF_X1 port map( D => n4220, CK => CLK, Q => 
                           REGISTERS_4_36_port, QN => n18059);
   REGISTERS_reg_4_35_inst : DFF_X1 port map( D => n4219, CK => CLK, Q => 
                           REGISTERS_4_35_port, QN => n18349);
   REGISTERS_reg_4_34_inst : DFF_X1 port map( D => n4218, CK => CLK, Q => 
                           REGISTERS_4_34_port, QN => n18060);
   REGISTERS_reg_4_33_inst : DFF_X1 port map( D => n4217, CK => CLK, Q => 
                           REGISTERS_4_33_port, QN => n18350);
   REGISTERS_reg_4_32_inst : DFF_X1 port map( D => n4216, CK => CLK, Q => 
                           REGISTERS_4_32_port, QN => n18351);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n4215, CK => CLK, Q => 
                           REGISTERS_4_31_port, QN => n18759);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n4214, CK => CLK, Q => 
                           REGISTERS_4_30_port, QN => n18352);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n4213, CK => CLK, Q => 
                           REGISTERS_4_29_port, QN => n18061);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n4212, CK => CLK, Q => 
                           REGISTERS_4_28_port, QN => n18353);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n4211, CK => CLK, Q => 
                           REGISTERS_4_27_port, QN => n17194);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n4210, CK => CLK, Q => 
                           REGISTERS_4_26_port, QN => n17810);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n4209, CK => CLK, Q => 
                           REGISTERS_4_25_port, QN => n17422);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n4208, CK => CLK, Q => 
                           REGISTERS_4_24_port, QN => n17423);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n4207, CK => CLK, Q => 
                           REGISTERS_4_23_port, QN => n17424);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n4206, CK => CLK, Q => 
                           REGISTERS_4_22_port, QN => n17195);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n4205, CK => CLK, Q => 
                           REGISTERS_4_21_port, QN => n17425);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n4204, CK => CLK, Q => 
                           REGISTERS_4_20_port, QN => n17811);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n4203, CK => CLK, Q => 
                           REGISTERS_4_19_port, QN => n17426);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n4202, CK => CLK, Q => 
                           REGISTERS_4_18_port, QN => n17196);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n4201, CK => CLK, Q => 
                           REGISTERS_4_17_port, QN => n17812);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n4200, CK => CLK, Q => 
                           REGISTERS_4_16_port, QN => n17197);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n4199, CK => CLK, Q => 
                           REGISTERS_4_15_port, QN => n18354);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n4198, CK => CLK, Q => 
                           REGISTERS_4_14_port, QN => n18355);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n4197, CK => CLK, Q => 
                           REGISTERS_4_13_port, QN => n18062);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n4196, CK => CLK, Q => 
                           REGISTERS_4_12_port, QN => n18356);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n4195, CK => CLK, Q => 
                           REGISTERS_4_11_port, QN => n18357);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n4194, CK => CLK, Q => 
                           REGISTERS_4_10_port, QN => n18358);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n4193, CK => CLK, Q => 
                           REGISTERS_4_9_port, QN => n18359);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n4192, CK => CLK, Q => 
                           REGISTERS_4_8_port, QN => n18360);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n4191, CK => CLK, Q => 
                           REGISTERS_4_7_port, QN => n18760);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n4190, CK => CLK, Q => 
                           REGISTERS_4_6_port, QN => n18761);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n4189, CK => CLK, Q => 
                           REGISTERS_4_5_port, QN => n18063);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n4188, CK => CLK, Q => 
                           REGISTERS_4_4_port, QN => n18064);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n4187, CK => CLK, Q => 
                           REGISTERS_4_3_port, QN => n18762);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n4186, CK => CLK, Q => 
                           REGISTERS_4_2_port, QN => n18361);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n4185, CK => CLK, Q => 
                           REGISTERS_4_1_port, QN => n18362);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n4184, CK => CLK, Q => 
                           REGISTERS_4_0_port, QN => n18363);
   REGISTERS_reg_5_63_inst : DFF_X1 port map( D => n4183, CK => CLK, Q => 
                           REGISTERS_5_63_port, QN => n16886);
   REGISTERS_reg_5_62_inst : DFF_X1 port map( D => n4182, CK => CLK, Q => 
                           REGISTERS_5_62_port, QN => n18364);
   REGISTERS_reg_5_61_inst : DFF_X1 port map( D => n4181, CK => CLK, Q => 
                           REGISTERS_5_61_port, QN => n18365);
   REGISTERS_reg_5_60_inst : DFF_X1 port map( D => n4180, CK => CLK, Q => 
                           REGISTERS_5_60_port, QN => n18366);
   REGISTERS_reg_5_59_inst : DFF_X1 port map( D => n4179, CK => CLK, Q => 
                           REGISTERS_5_59_port, QN => n18367);
   REGISTERS_reg_5_58_inst : DFF_X1 port map( D => n4178, CK => CLK, Q => 
                           REGISTERS_5_58_port, QN => n18763);
   REGISTERS_reg_5_57_inst : DFF_X1 port map( D => n4177, CK => CLK, Q => 
                           REGISTERS_5_57_port, QN => n18368);
   REGISTERS_reg_5_56_inst : DFF_X1 port map( D => n4176, CK => CLK, Q => 
                           REGISTERS_5_56_port, QN => n18764);
   REGISTERS_reg_5_55_inst : DFF_X1 port map( D => n4175, CK => CLK, Q => 
                           REGISTERS_5_55_port, QN => n18765);
   REGISTERS_reg_5_54_inst : DFF_X1 port map( D => n4174, CK => CLK, Q => 
                           REGISTERS_5_54_port, QN => n18766);
   REGISTERS_reg_5_53_inst : DFF_X1 port map( D => n4173, CK => CLK, Q => 
                           REGISTERS_5_53_port, QN => n18369);
   REGISTERS_reg_5_52_inst : DFF_X1 port map( D => n4172, CK => CLK, Q => 
                           REGISTERS_5_52_port, QN => n18767);
   REGISTERS_reg_5_51_inst : DFF_X1 port map( D => n4171, CK => CLK, Q => 
                           REGISTERS_5_51_port, QN => n18065);
   REGISTERS_reg_5_50_inst : DFF_X1 port map( D => n4170, CK => CLK, Q => 
                           REGISTERS_5_50_port, QN => n18768);
   REGISTERS_reg_5_49_inst : DFF_X1 port map( D => n4169, CK => CLK, Q => 
                           REGISTERS_5_49_port, QN => n18370);
   REGISTERS_reg_5_48_inst : DFF_X1 port map( D => n4168, CK => CLK, Q => 
                           REGISTERS_5_48_port, QN => n18371);
   REGISTERS_reg_5_47_inst : DFF_X1 port map( D => n4167, CK => CLK, Q => 
                           REGISTERS_5_47_port, QN => n18769);
   REGISTERS_reg_5_46_inst : DFF_X1 port map( D => n4166, CK => CLK, Q => 
                           REGISTERS_5_46_port, QN => n18770);
   REGISTERS_reg_5_45_inst : DFF_X1 port map( D => n4165, CK => CLK, Q => 
                           REGISTERS_5_45_port, QN => n18372);
   REGISTERS_reg_5_44_inst : DFF_X1 port map( D => n4164, CK => CLK, Q => 
                           REGISTERS_5_44_port, QN => n18373);
   REGISTERS_reg_5_43_inst : DFF_X1 port map( D => n4163, CK => CLK, Q => 
                           REGISTERS_5_43_port, QN => n18374);
   REGISTERS_reg_5_42_inst : DFF_X1 port map( D => n4162, CK => CLK, Q => 
                           REGISTERS_5_42_port, QN => n18771);
   REGISTERS_reg_5_41_inst : DFF_X1 port map( D => n4161, CK => CLK, Q => 
                           REGISTERS_5_41_port, QN => n18772);
   REGISTERS_reg_5_40_inst : DFF_X1 port map( D => n4160, CK => CLK, Q => 
                           REGISTERS_5_40_port, QN => n18773);
   REGISTERS_reg_5_39_inst : DFF_X1 port map( D => n4159, CK => CLK, Q => 
                           REGISTERS_5_39_port, QN => n18774);
   REGISTERS_reg_5_38_inst : DFF_X1 port map( D => n4158, CK => CLK, Q => 
                           REGISTERS_5_38_port, QN => n18775);
   REGISTERS_reg_5_37_inst : DFF_X1 port map( D => n4157, CK => CLK, Q => 
                           REGISTERS_5_37_port, QN => n18375);
   REGISTERS_reg_5_36_inst : DFF_X1 port map( D => n4156, CK => CLK, Q => 
                           REGISTERS_5_36_port, QN => n18776);
   REGISTERS_reg_5_35_inst : DFF_X1 port map( D => n4155, CK => CLK, Q => 
                           REGISTERS_5_35_port, QN => n18777);
   REGISTERS_reg_5_34_inst : DFF_X1 port map( D => n4154, CK => CLK, Q => 
                           REGISTERS_5_34_port, QN => n18376);
   REGISTERS_reg_5_33_inst : DFF_X1 port map( D => n4153, CK => CLK, Q => 
                           REGISTERS_5_33_port, QN => n18778);
   REGISTERS_reg_5_32_inst : DFF_X1 port map( D => n4152, CK => CLK, Q => 
                           REGISTERS_5_32_port, QN => n18779);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n4151, CK => CLK, Q => 
                           REGISTERS_5_31_port, QN => n18780);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n4150, CK => CLK, Q => 
                           REGISTERS_5_30_port, QN => n18377);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n4149, CK => CLK, Q => 
                           REGISTERS_5_29_port, QN => n18378);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n4148, CK => CLK, Q => 
                           REGISTERS_5_28_port, QN => n18379);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n4147, CK => CLK, Q => 
                           REGISTERS_5_27_port, QN => n17427);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n4146, CK => CLK, Q => 
                           REGISTERS_5_26_port, QN => n17428);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n4145, CK => CLK, Q => 
                           REGISTERS_5_25_port, QN => n17429);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n4144, CK => CLK, Q => 
                           REGISTERS_5_24_port, QN => n17430);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n4143, CK => CLK, Q => 
                           REGISTERS_5_23_port, QN => n17198);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n4142, CK => CLK, Q => 
                           REGISTERS_5_22_port, QN => n17813);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n4141, CK => CLK, Q => 
                           REGISTERS_5_21_port, QN => n17814);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n4140, CK => CLK, Q => 
                           REGISTERS_5_20_port, QN => n17815);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n4139, CK => CLK, Q => 
                           REGISTERS_5_19_port, QN => n17816);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n4138, CK => CLK, Q => 
                           REGISTERS_5_18_port, QN => n17431);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n4137, CK => CLK, Q => 
                           REGISTERS_5_17_port, QN => n17199);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n4136, CK => n13730, Q => 
                           REGISTERS_5_16_port, QN => n17817);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n4135, CK => CLK, Q => 
                           REGISTERS_5_15_port, QN => n18066);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n4134, CK => CLK, Q => 
                           REGISTERS_5_14_port, QN => n18781);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n4133, CK => CLK, Q => 
                           REGISTERS_5_13_port, QN => n18067);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n4132, CK => CLK, Q => 
                           REGISTERS_5_12_port, QN => n18380);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n4131, CK => CLK, Q => 
                           REGISTERS_5_11_port, QN => n18068);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n4130, CK => CLK, Q => 
                           REGISTERS_5_10_port, QN => n18782);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n4129, CK => CLK, Q => 
                           REGISTERS_5_9_port, QN => n18783);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n4128, CK => CLK, Q => 
                           REGISTERS_5_8_port, QN => n18784);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n4127, CK => CLK, Q => 
                           REGISTERS_5_7_port, QN => n18069);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n4126, CK => CLK, Q => 
                           REGISTERS_5_6_port, QN => n18381);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n4125, CK => CLK, Q => 
                           REGISTERS_5_5_port, QN => n18382);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n4124, CK => CLK, Q => 
                           REGISTERS_5_4_port, QN => n18383);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n4123, CK => CLK, Q => 
                           REGISTERS_5_3_port, QN => n18384);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n4122, CK => CLK, Q => 
                           REGISTERS_5_2_port, QN => n18385);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n4121, CK => CLK, Q => 
                           REGISTERS_5_1_port, QN => n18386);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n4120, CK => CLK, Q => 
                           REGISTERS_5_0_port, QN => n18387);
   REGISTERS_reg_6_63_inst : DFF_X1 port map( D => n4119, CK => CLK, Q => 
                           REGISTERS_6_63_port, QN => n16964);
   REGISTERS_reg_6_62_inst : DFF_X1 port map( D => n4118, CK => CLK, Q => 
                           REGISTERS_6_62_port, QN => n18388);
   REGISTERS_reg_6_61_inst : DFF_X1 port map( D => n4117, CK => CLK, Q => 
                           REGISTERS_6_61_port, QN => n18785);
   REGISTERS_reg_6_60_inst : DFF_X1 port map( D => n4116, CK => CLK, Q => 
                           REGISTERS_6_60_port, QN => n18389);
   REGISTERS_reg_6_59_inst : DFF_X1 port map( D => n4115, CK => CLK, Q => 
                           REGISTERS_6_59_port, QN => n18390);
   REGISTERS_reg_6_58_inst : DFF_X1 port map( D => n4114, CK => CLK, Q => 
                           REGISTERS_6_58_port, QN => n18391);
   REGISTERS_reg_6_57_inst : DFF_X1 port map( D => n4113, CK => CLK, Q => 
                           REGISTERS_6_57_port, QN => n18392);
   REGISTERS_reg_6_56_inst : DFF_X1 port map( D => n4112, CK => CLK, Q => 
                           REGISTERS_6_56_port, QN => n18786);
   REGISTERS_reg_6_55_inst : DFF_X1 port map( D => n4111, CK => CLK, Q => 
                           REGISTERS_6_55_port, QN => n18393);
   REGISTERS_reg_6_54_inst : DFF_X1 port map( D => n4110, CK => CLK, Q => 
                           REGISTERS_6_54_port, QN => n18070);
   REGISTERS_reg_6_53_inst : DFF_X1 port map( D => n4109, CK => CLK, Q => 
                           REGISTERS_6_53_port, QN => n18394);
   REGISTERS_reg_6_52_inst : DFF_X1 port map( D => n4108, CK => CLK, Q => 
                           REGISTERS_6_52_port, QN => n18071);
   REGISTERS_reg_6_51_inst : DFF_X1 port map( D => n4107, CK => CLK, Q => 
                           REGISTERS_6_51_port, QN => n18395);
   REGISTERS_reg_6_50_inst : DFF_X1 port map( D => n4106, CK => CLK, Q => 
                           REGISTERS_6_50_port, QN => n18396);
   REGISTERS_reg_6_49_inst : DFF_X1 port map( D => n4105, CK => CLK, Q => 
                           REGISTERS_6_49_port, QN => n18787);
   REGISTERS_reg_6_48_inst : DFF_X1 port map( D => n4104, CK => CLK, Q => 
                           REGISTERS_6_48_port, QN => n18788);
   REGISTERS_reg_6_47_inst : DFF_X1 port map( D => n4103, CK => CLK, Q => 
                           REGISTERS_6_47_port, QN => n18072);
   REGISTERS_reg_6_46_inst : DFF_X1 port map( D => n4102, CK => CLK, Q => 
                           REGISTERS_6_46_port, QN => n18397);
   REGISTERS_reg_6_45_inst : DFF_X1 port map( D => n4101, CK => CLK, Q => 
                           REGISTERS_6_45_port, QN => n18398);
   REGISTERS_reg_6_44_inst : DFF_X1 port map( D => n4100, CK => CLK, Q => 
                           REGISTERS_6_44_port, QN => n18073);
   REGISTERS_reg_6_43_inst : DFF_X1 port map( D => n4099, CK => CLK, Q => 
                           REGISTERS_6_43_port, QN => n18789);
   REGISTERS_reg_6_42_inst : DFF_X1 port map( D => n4098, CK => CLK, Q => 
                           REGISTERS_6_42_port, QN => n18399);
   REGISTERS_reg_6_41_inst : DFF_X1 port map( D => n4097, CK => CLK, Q => 
                           REGISTERS_6_41_port, QN => n18400);
   REGISTERS_reg_6_40_inst : DFF_X1 port map( D => n4096, CK => CLK, Q => 
                           REGISTERS_6_40_port, QN => n18790);
   REGISTERS_reg_6_39_inst : DFF_X1 port map( D => n4095, CK => CLK, Q => 
                           REGISTERS_6_39_port, QN => n18074);
   REGISTERS_reg_6_38_inst : DFF_X1 port map( D => n4094, CK => CLK, Q => 
                           REGISTERS_6_38_port, QN => n18075);
   REGISTERS_reg_6_37_inst : DFF_X1 port map( D => n4093, CK => CLK, Q => 
                           REGISTERS_6_37_port, QN => n18791);
   REGISTERS_reg_6_36_inst : DFF_X1 port map( D => n4092, CK => CLK, Q => 
                           REGISTERS_6_36_port, QN => n18076);
   REGISTERS_reg_6_35_inst : DFF_X1 port map( D => n4091, CK => CLK, Q => 
                           REGISTERS_6_35_port, QN => n18077);
   REGISTERS_reg_6_34_inst : DFF_X1 port map( D => n4090, CK => CLK, Q => 
                           REGISTERS_6_34_port, QN => n18401);
   REGISTERS_reg_6_33_inst : DFF_X1 port map( D => n4089, CK => CLK, Q => 
                           REGISTERS_6_33_port, QN => n18402);
   REGISTERS_reg_6_32_inst : DFF_X1 port map( D => n4088, CK => CLK, Q => 
                           REGISTERS_6_32_port, QN => n18078);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n4087, CK => CLK, Q => 
                           REGISTERS_6_31_port, QN => n18079);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n4086, CK => CLK, Q => 
                           REGISTERS_6_30_port, QN => n18403);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n4085, CK => CLK, Q => 
                           REGISTERS_6_29_port, QN => n18404);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n4084, CK => CLK, Q => 
                           REGISTERS_6_28_port, QN => n18405);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n4083, CK => CLK, Q => 
                           REGISTERS_6_27_port, QN => n17432);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n4082, CK => CLK, Q => 
                           REGISTERS_6_26_port, QN => n17200);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n4081, CK => CLK, Q => 
                           REGISTERS_6_25_port, QN => n17818);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n4080, CK => CLK, Q => 
                           REGISTERS_6_24_port, QN => n17433);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n4079, CK => CLK, Q => 
                           REGISTERS_6_23_port, QN => n17819);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n4078, CK => CLK, Q => 
                           REGISTERS_6_22_port, QN => n17434);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n4077, CK => CLK, Q => 
                           REGISTERS_6_21_port, QN => n17435);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n4076, CK => CLK, Q => 
                           REGISTERS_6_20_port, QN => n17436);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n4075, CK => CLK, Q => 
                           REGISTERS_6_19_port, QN => n17201);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n4074, CK => CLK, Q => 
                           REGISTERS_6_18_port, QN => n17437);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n4073, CK => CLK, Q => 
                           REGISTERS_6_17_port, QN => n17202);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n4072, CK => CLK, Q => 
                           REGISTERS_6_16_port, QN => n17203);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n4071, CK => CLK, Q => 
                           REGISTERS_6_15_port, QN => n18406);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n4070, CK => CLK, Q => 
                           REGISTERS_6_14_port, QN => n18407);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n4069, CK => CLK, Q => 
                           REGISTERS_6_13_port, QN => n18792);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n4068, CK => CLK, Q => 
                           REGISTERS_6_12_port, QN => n18408);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n4067, CK => CLK, Q => 
                           REGISTERS_6_11_port, QN => n18409);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n4066, CK => CLK, Q => 
                           REGISTERS_6_10_port, QN => n18410);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n4065, CK => CLK, Q => 
                           REGISTERS_6_9_port, QN => n18411);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n4064, CK => CLK, Q => 
                           REGISTERS_6_8_port, QN => n18080);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n4063, CK => CLK, Q => 
                           REGISTERS_6_7_port, QN => n18793);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n4062, CK => CLK, Q => 
                           REGISTERS_6_6_port, QN => n18412);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n4061, CK => CLK, Q => 
                           REGISTERS_6_5_port, QN => n18413);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n4060, CK => CLK, Q => 
                           REGISTERS_6_4_port, QN => n18414);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n4059, CK => CLK, Q => 
                           REGISTERS_6_3_port, QN => n18081);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n4058, CK => CLK, Q => 
                           REGISTERS_6_2_port, QN => n18415);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n4057, CK => CLK, Q => 
                           REGISTERS_6_1_port, QN => n18794);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n4056, CK => CLK, Q => 
                           REGISTERS_6_0_port, QN => n18795);
   REGISTERS_reg_7_63_inst : DFF_X1 port map( D => n4055, CK => CLK, Q => 
                           REGISTERS_7_63_port, QN => n17107);
   REGISTERS_reg_7_62_inst : DFF_X1 port map( D => n4054, CK => CLK, Q => 
                           REGISTERS_7_62_port, QN => n18416);
   REGISTERS_reg_7_61_inst : DFF_X1 port map( D => n4053, CK => CLK, Q => 
                           REGISTERS_7_61_port, QN => n18417);
   REGISTERS_reg_7_60_inst : DFF_X1 port map( D => n4052, CK => CLK, Q => 
                           REGISTERS_7_60_port, QN => n18418);
   REGISTERS_reg_7_59_inst : DFF_X1 port map( D => n4051, CK => CLK, Q => 
                           REGISTERS_7_59_port, QN => n18082);
   REGISTERS_reg_7_58_inst : DFF_X1 port map( D => n4050, CK => CLK, Q => 
                           REGISTERS_7_58_port, QN => n18083);
   REGISTERS_reg_7_57_inst : DFF_X1 port map( D => n4049, CK => CLK, Q => 
                           REGISTERS_7_57_port, QN => n18419);
   REGISTERS_reg_7_56_inst : DFF_X1 port map( D => n4048, CK => CLK, Q => 
                           REGISTERS_7_56_port, QN => n18420);
   REGISTERS_reg_7_55_inst : DFF_X1 port map( D => n4047, CK => CLK, Q => 
                           REGISTERS_7_55_port, QN => n18421);
   REGISTERS_reg_7_54_inst : DFF_X1 port map( D => n4046, CK => CLK, Q => 
                           REGISTERS_7_54_port, QN => n18084);
   REGISTERS_reg_7_53_inst : DFF_X1 port map( D => n4045, CK => CLK, Q => 
                           REGISTERS_7_53_port, QN => n18085);
   REGISTERS_reg_7_52_inst : DFF_X1 port map( D => n4044, CK => CLK, Q => 
                           REGISTERS_7_52_port, QN => n18422);
   REGISTERS_reg_7_51_inst : DFF_X1 port map( D => n4043, CK => CLK, Q => 
                           REGISTERS_7_51_port, QN => n18796);
   REGISTERS_reg_7_50_inst : DFF_X1 port map( D => n4042, CK => CLK, Q => 
                           REGISTERS_7_50_port, QN => n18086);
   REGISTERS_reg_7_49_inst : DFF_X1 port map( D => n4041, CK => CLK, Q => 
                           REGISTERS_7_49_port, QN => n18423);
   REGISTERS_reg_7_48_inst : DFF_X1 port map( D => n4040, CK => CLK, Q => 
                           REGISTERS_7_48_port, QN => n18087);
   REGISTERS_reg_7_47_inst : DFF_X1 port map( D => n4039, CK => CLK, Q => 
                           REGISTERS_7_47_port, QN => n18088);
   REGISTERS_reg_7_46_inst : DFF_X1 port map( D => n4038, CK => CLK, Q => 
                           REGISTERS_7_46_port, QN => n18424);
   REGISTERS_reg_7_45_inst : DFF_X1 port map( D => n4037, CK => CLK, Q => 
                           REGISTERS_7_45_port, QN => n18089);
   REGISTERS_reg_7_44_inst : DFF_X1 port map( D => n4036, CK => CLK, Q => 
                           REGISTERS_7_44_port, QN => n18797);
   REGISTERS_reg_7_43_inst : DFF_X1 port map( D => n4035, CK => CLK, Q => 
                           REGISTERS_7_43_port, QN => n18090);
   REGISTERS_reg_7_42_inst : DFF_X1 port map( D => n4034, CK => CLK, Q => 
                           REGISTERS_7_42_port, QN => n18425);
   REGISTERS_reg_7_41_inst : DFF_X1 port map( D => n4033, CK => CLK, Q => 
                           REGISTERS_7_41_port, QN => n18426);
   REGISTERS_reg_7_40_inst : DFF_X1 port map( D => n4032, CK => CLK, Q => 
                           REGISTERS_7_40_port, QN => n18427);
   REGISTERS_reg_7_39_inst : DFF_X1 port map( D => n4031, CK => CLK, Q => 
                           REGISTERS_7_39_port, QN => n18428);
   REGISTERS_reg_7_38_inst : DFF_X1 port map( D => n4030, CK => CLK, Q => 
                           REGISTERS_7_38_port, QN => n18091);
   REGISTERS_reg_7_37_inst : DFF_X1 port map( D => n4029, CK => CLK, Q => 
                           REGISTERS_7_37_port, QN => n18092);
   REGISTERS_reg_7_36_inst : DFF_X1 port map( D => n4028, CK => CLK, Q => 
                           REGISTERS_7_36_port, QN => n18429);
   REGISTERS_reg_7_35_inst : DFF_X1 port map( D => n4027, CK => CLK, Q => 
                           REGISTERS_7_35_port, QN => n18093);
   REGISTERS_reg_7_34_inst : DFF_X1 port map( D => n4026, CK => CLK, Q => 
                           REGISTERS_7_34_port, QN => n18430);
   REGISTERS_reg_7_33_inst : DFF_X1 port map( D => n4025, CK => CLK, Q => 
                           REGISTERS_7_33_port, QN => n18431);
   REGISTERS_reg_7_32_inst : DFF_X1 port map( D => n4024, CK => CLK, Q => 
                           REGISTERS_7_32_port, QN => n18432);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n4023, CK => CLK, Q => 
                           REGISTERS_7_31_port, QN => n18433);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n4022, CK => CLK, Q => 
                           REGISTERS_7_30_port, QN => n18094);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n4021, CK => CLK, Q => 
                           REGISTERS_7_29_port, QN => n18434);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n4020, CK => CLK, Q => 
                           REGISTERS_7_28_port, QN => n18095);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n4019, CK => CLK, Q => 
                           REGISTERS_7_27_port, QN => n17438);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n4018, CK => CLK, Q => 
                           REGISTERS_7_26_port, QN => n17204);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n4017, CK => CLK, Q => 
                           REGISTERS_7_25_port, QN => n17205);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n4016, CK => CLK, Q => 
                           REGISTERS_7_24_port, QN => n17206);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n4015, CK => CLK, Q => 
                           REGISTERS_7_23_port, QN => n17207);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n4014, CK => CLK, Q => 
                           REGISTERS_7_22_port, QN => n17439);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n4013, CK => CLK, Q => 
                           REGISTERS_7_21_port, QN => n17208);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n4012, CK => CLK, Q => 
                           REGISTERS_7_20_port, QN => n17440);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n4011, CK => CLK, Q => 
                           REGISTERS_7_19_port, QN => n17441);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n4010, CK => CLK, Q => 
                           REGISTERS_7_18_port, QN => n17209);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n4009, CK => CLK, Q => 
                           REGISTERS_7_17_port, QN => n17442);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n4008, CK => CLK, Q => 
                           REGISTERS_7_16_port, QN => n17443);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n4007, CK => CLK, Q => 
                           REGISTERS_7_15_port, QN => n18435);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n4006, CK => CLK, Q => 
                           REGISTERS_7_14_port, QN => n18096);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n4005, CK => CLK, Q => 
                           REGISTERS_7_13_port, QN => n18798);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n4004, CK => CLK, Q => 
                           REGISTERS_7_12_port, QN => n18097);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n4003, CK => CLK, Q => 
                           REGISTERS_7_11_port, QN => n18098);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n4002, CK => CLK, Q => 
                           REGISTERS_7_10_port, QN => n18799);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n4001, CK => CLK, Q => 
                           REGISTERS_7_9_port, QN => n18436);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n4000, CK => CLK, Q => 
                           REGISTERS_7_8_port, QN => n18437);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n3999, CK => CLK, Q => 
                           REGISTERS_7_7_port, QN => n18438);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n3998, CK => CLK, Q => 
                           REGISTERS_7_6_port, QN => n18439);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n3997, CK => CLK, Q => 
                           REGISTERS_7_5_port, QN => n18440);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n3996, CK => CLK, Q => 
                           REGISTERS_7_4_port, QN => n18099);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n3995, CK => CLK, Q => 
                           REGISTERS_7_3_port, QN => n18100);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n3994, CK => CLK, Q => 
                           REGISTERS_7_2_port, QN => n18101);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n3993, CK => CLK, Q => 
                           REGISTERS_7_1_port, QN => n18102);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n3992, CK => CLK, Q => 
                           REGISTERS_7_0_port, QN => n18103);
   REGISTERS_reg_8_63_inst : DFF_X1 port map( D => n3991, CK => CLK, Q => 
                           REGISTERS_8_63_port, QN => n16883);
   REGISTERS_reg_8_62_inst : DFF_X1 port map( D => n3990, CK => CLK, Q => 
                           REGISTERS_8_62_port, QN => n18441);
   REGISTERS_reg_8_61_inst : DFF_X1 port map( D => n3989, CK => CLK, Q => 
                           REGISTERS_8_61_port, QN => n18442);
   REGISTERS_reg_8_60_inst : DFF_X1 port map( D => n3988, CK => CLK, Q => 
                           REGISTERS_8_60_port, QN => n18800);
   REGISTERS_reg_8_59_inst : DFF_X1 port map( D => n3987, CK => CLK, Q => 
                           REGISTERS_8_59_port, QN => n18104);
   REGISTERS_reg_8_58_inst : DFF_X1 port map( D => n3986, CK => CLK, Q => 
                           REGISTERS_8_58_port, QN => n18443);
   REGISTERS_reg_8_57_inst : DFF_X1 port map( D => n3985, CK => CLK, Q => 
                           REGISTERS_8_57_port, QN => n18444);
   REGISTERS_reg_8_56_inst : DFF_X1 port map( D => n3984, CK => CLK, Q => 
                           REGISTERS_8_56_port, QN => n18445);
   REGISTERS_reg_8_55_inst : DFF_X1 port map( D => n3983, CK => CLK, Q => 
                           REGISTERS_8_55_port, QN => n18105);
   REGISTERS_reg_8_54_inst : DFF_X1 port map( D => n3982, CK => CLK, Q => 
                           REGISTERS_8_54_port, QN => n18446);
   REGISTERS_reg_8_53_inst : DFF_X1 port map( D => n3981, CK => CLK, Q => 
                           REGISTERS_8_53_port, QN => n18447);
   REGISTERS_reg_8_52_inst : DFF_X1 port map( D => n3980, CK => CLK, Q => 
                           REGISTERS_8_52_port, QN => n18106);
   REGISTERS_reg_8_51_inst : DFF_X1 port map( D => n3979, CK => CLK, Q => 
                           REGISTERS_8_51_port, QN => n18448);
   REGISTERS_reg_8_50_inst : DFF_X1 port map( D => n3978, CK => n13730, Q => 
                           REGISTERS_8_50_port, QN => n18449);
   REGISTERS_reg_8_49_inst : DFF_X1 port map( D => n3977, CK => CLK, Q => 
                           REGISTERS_8_49_port, QN => n18450);
   REGISTERS_reg_8_48_inst : DFF_X1 port map( D => n3976, CK => CLK, Q => 
                           REGISTERS_8_48_port, QN => n18451);
   REGISTERS_reg_8_47_inst : DFF_X1 port map( D => n3975, CK => CLK, Q => 
                           REGISTERS_8_47_port, QN => n18452);
   REGISTERS_reg_8_46_inst : DFF_X1 port map( D => n3974, CK => CLK, Q => 
                           REGISTERS_8_46_port, QN => n18453);
   REGISTERS_reg_8_45_inst : DFF_X1 port map( D => n3973, CK => CLK, Q => 
                           REGISTERS_8_45_port, QN => n18454);
   REGISTERS_reg_8_44_inst : DFF_X1 port map( D => n3972, CK => CLK, Q => 
                           REGISTERS_8_44_port, QN => n18801);
   REGISTERS_reg_8_43_inst : DFF_X1 port map( D => n3971, CK => CLK, Q => 
                           REGISTERS_8_43_port, QN => n18107);
   REGISTERS_reg_8_42_inst : DFF_X1 port map( D => n3970, CK => CLK, Q => 
                           REGISTERS_8_42_port, QN => n18802);
   REGISTERS_reg_8_41_inst : DFF_X1 port map( D => n3969, CK => CLK, Q => 
                           REGISTERS_8_41_port, QN => n18455);
   REGISTERS_reg_8_40_inst : DFF_X1 port map( D => n3968, CK => CLK, Q => 
                           REGISTERS_8_40_port, QN => n18108);
   REGISTERS_reg_8_39_inst : DFF_X1 port map( D => n3967, CK => CLK, Q => 
                           REGISTERS_8_39_port, QN => n18456);
   REGISTERS_reg_8_38_inst : DFF_X1 port map( D => n3966, CK => CLK, Q => 
                           REGISTERS_8_38_port, QN => n18457);
   REGISTERS_reg_8_37_inst : DFF_X1 port map( D => n3965, CK => CLK, Q => 
                           REGISTERS_8_37_port, QN => n18109);
   REGISTERS_reg_8_36_inst : DFF_X1 port map( D => n3964, CK => CLK, Q => 
                           REGISTERS_8_36_port, QN => n18458);
   REGISTERS_reg_8_35_inst : DFF_X1 port map( D => n3963, CK => CLK, Q => 
                           REGISTERS_8_35_port, QN => n18110);
   REGISTERS_reg_8_34_inst : DFF_X1 port map( D => n3962, CK => CLK, Q => 
                           REGISTERS_8_34_port, QN => n18459);
   REGISTERS_reg_8_33_inst : DFF_X1 port map( D => n3961, CK => CLK, Q => 
                           REGISTERS_8_33_port, QN => n18111);
   REGISTERS_reg_8_32_inst : DFF_X1 port map( D => n3960, CK => CLK, Q => 
                           REGISTERS_8_32_port, QN => n18112);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n3959, CK => CLK, Q => 
                           REGISTERS_8_31_port, QN => n18113);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n3958, CK => CLK, Q => 
                           REGISTERS_8_30_port, QN => n18460);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n3957, CK => CLK, Q => 
                           REGISTERS_8_29_port, QN => n18461);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n3956, CK => CLK, Q => 
                           REGISTERS_8_28_port, QN => n18114);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n3955, CK => CLK, Q => 
                           REGISTERS_8_27_port, QN => n17820);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n3954, CK => CLK, Q => 
                           REGISTERS_8_26_port, QN => n17821);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n3953, CK => CLK, Q => 
                           REGISTERS_8_25_port, QN => n17444);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n3952, CK => CLK, Q => 
                           REGISTERS_8_24_port, QN => n17445);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n3951, CK => CLK, Q => 
                           REGISTERS_8_23_port, QN => n17446);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n3950, CK => CLK, Q => 
                           REGISTERS_8_22_port, QN => n17447);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n3949, CK => CLK, Q => 
                           REGISTERS_8_21_port, QN => n17210);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n3948, CK => CLK, Q => 
                           REGISTERS_8_20_port, QN => n17448);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n3947, CK => CLK, Q => 
                           REGISTERS_8_19_port, QN => n17211);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n3946, CK => CLK, Q => 
                           REGISTERS_8_18_port, QN => n17822);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n3945, CK => CLK, Q => 
                           REGISTERS_8_17_port, QN => n17449);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n3944, CK => CLK, Q => 
                           REGISTERS_8_16_port, QN => n17450);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n3943, CK => CLK, Q => 
                           REGISTERS_8_15_port, QN => n18462);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n3942, CK => CLK, Q => 
                           REGISTERS_8_14_port, QN => n18803);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n3941, CK => CLK, Q => 
                           REGISTERS_8_13_port, QN => n18115);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n3940, CK => CLK, Q => 
                           REGISTERS_8_12_port, QN => n18463);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n3939, CK => CLK, Q => 
                           REGISTERS_8_11_port, QN => n18464);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n3938, CK => CLK, Q => 
                           REGISTERS_8_10_port, QN => n18116);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n3937, CK => CLK, Q => 
                           REGISTERS_8_9_port, QN => n18465);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n3936, CK => CLK, Q => 
                           REGISTERS_8_8_port, QN => n18466);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n3935, CK => CLK, Q => 
                           REGISTERS_8_7_port, QN => n18117);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n3934, CK => CLK, Q => 
                           REGISTERS_8_6_port, QN => n18467);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n3933, CK => CLK, Q => 
                           REGISTERS_8_5_port, QN => n18468);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n3932, CK => CLK, Q => 
                           REGISTERS_8_4_port, QN => n18118);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n3931, CK => CLK, Q => 
                           REGISTERS_8_3_port, QN => n18469);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n3930, CK => CLK, Q => 
                           REGISTERS_8_2_port, QN => n18119);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n3929, CK => CLK, Q => 
                           REGISTERS_8_1_port, QN => n18470);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n3928, CK => CLK, Q => 
                           REGISTERS_8_0_port, QN => n18471);
   REGISTERS_reg_9_63_inst : DFF_X1 port map( D => n3927, CK => CLK, Q => 
                           REGISTERS_9_63_port, QN => n16887);
   REGISTERS_reg_9_62_inst : DFF_X1 port map( D => n3926, CK => CLK, Q => 
                           REGISTERS_9_62_port, QN => n18120);
   REGISTERS_reg_9_61_inst : DFF_X1 port map( D => n3925, CK => CLK, Q => 
                           REGISTERS_9_61_port, QN => n18804);
   REGISTERS_reg_9_60_inst : DFF_X1 port map( D => n3924, CK => CLK, Q => 
                           REGISTERS_9_60_port, QN => n18805);
   REGISTERS_reg_9_59_inst : DFF_X1 port map( D => n3923, CK => CLK, Q => 
                           REGISTERS_9_59_port, QN => n18121);
   REGISTERS_reg_9_58_inst : DFF_X1 port map( D => n3922, CK => CLK, Q => 
                           REGISTERS_9_58_port, QN => n18122);
   REGISTERS_reg_9_57_inst : DFF_X1 port map( D => n3921, CK => CLK, Q => 
                           REGISTERS_9_57_port, QN => n18472);
   REGISTERS_reg_9_56_inst : DFF_X1 port map( D => n3920, CK => CLK, Q => 
                           REGISTERS_9_56_port, QN => n18123);
   REGISTERS_reg_9_55_inst : DFF_X1 port map( D => n3919, CK => CLK, Q => 
                           REGISTERS_9_55_port, QN => n18473);
   REGISTERS_reg_9_54_inst : DFF_X1 port map( D => n3918, CK => CLK, Q => 
                           REGISTERS_9_54_port, QN => n18474);
   REGISTERS_reg_9_53_inst : DFF_X1 port map( D => n3917, CK => CLK, Q => 
                           REGISTERS_9_53_port, QN => n18475);
   REGISTERS_reg_9_52_inst : DFF_X1 port map( D => n3916, CK => CLK, Q => 
                           REGISTERS_9_52_port, QN => n18806);
   REGISTERS_reg_9_51_inst : DFF_X1 port map( D => n3915, CK => CLK, Q => 
                           REGISTERS_9_51_port, QN => n18124);
   REGISTERS_reg_9_50_inst : DFF_X1 port map( D => n3914, CK => CLK, Q => 
                           REGISTERS_9_50_port, QN => n18125);
   REGISTERS_reg_9_49_inst : DFF_X1 port map( D => n3913, CK => CLK, Q => 
                           REGISTERS_9_49_port, QN => n18476);
   REGISTERS_reg_9_48_inst : DFF_X1 port map( D => n3912, CK => CLK, Q => 
                           REGISTERS_9_48_port, QN => n18126);
   REGISTERS_reg_9_47_inst : DFF_X1 port map( D => n3911, CK => CLK, Q => 
                           REGISTERS_9_47_port, QN => n18127);
   REGISTERS_reg_9_46_inst : DFF_X1 port map( D => n3910, CK => CLK, Q => 
                           REGISTERS_9_46_port, QN => n18477);
   REGISTERS_reg_9_45_inst : DFF_X1 port map( D => n3909, CK => CLK, Q => 
                           REGISTERS_9_45_port, QN => n18478);
   REGISTERS_reg_9_44_inst : DFF_X1 port map( D => n3908, CK => CLK, Q => 
                           REGISTERS_9_44_port, QN => n18479);
   REGISTERS_reg_9_43_inst : DFF_X1 port map( D => n3907, CK => CLK, Q => 
                           REGISTERS_9_43_port, QN => n18480);
   REGISTERS_reg_9_42_inst : DFF_X1 port map( D => n3906, CK => CLK, Q => 
                           REGISTERS_9_42_port, QN => n18128);
   REGISTERS_reg_9_41_inst : DFF_X1 port map( D => n3905, CK => CLK, Q => 
                           REGISTERS_9_41_port, QN => n18481);
   REGISTERS_reg_9_40_inst : DFF_X1 port map( D => n3904, CK => CLK, Q => 
                           REGISTERS_9_40_port, QN => n18482);
   REGISTERS_reg_9_39_inst : DFF_X1 port map( D => n3903, CK => CLK, Q => 
                           REGISTERS_9_39_port, QN => n18483);
   REGISTERS_reg_9_38_inst : DFF_X1 port map( D => n3902, CK => CLK, Q => 
                           REGISTERS_9_38_port, QN => n18129);
   REGISTERS_reg_9_37_inst : DFF_X1 port map( D => n3901, CK => CLK, Q => 
                           REGISTERS_9_37_port, QN => n18484);
   REGISTERS_reg_9_36_inst : DFF_X1 port map( D => n3900, CK => CLK, Q => 
                           REGISTERS_9_36_port, QN => n18485);
   REGISTERS_reg_9_35_inst : DFF_X1 port map( D => n3899, CK => CLK, Q => 
                           REGISTERS_9_35_port, QN => n18130);
   REGISTERS_reg_9_34_inst : DFF_X1 port map( D => n3898, CK => CLK, Q => 
                           REGISTERS_9_34_port, QN => n18486);
   REGISTERS_reg_9_33_inst : DFF_X1 port map( D => n3897, CK => CLK, Q => 
                           REGISTERS_9_33_port, QN => n18487);
   REGISTERS_reg_9_32_inst : DFF_X1 port map( D => n3896, CK => CLK, Q => 
                           REGISTERS_9_32_port, QN => n18488);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n3895, CK => CLK, Q => 
                           REGISTERS_9_31_port, QN => n18489);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n3894, CK => CLK, Q => 
                           REGISTERS_9_30_port, QN => n18131);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n3893, CK => CLK, Q => 
                           REGISTERS_9_29_port, QN => n18132);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n3892, CK => CLK, Q => 
                           REGISTERS_9_28_port, QN => n18490);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n3891, CK => CLK, Q => 
                           REGISTERS_9_27_port, QN => n17823);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n3890, CK => CLK, Q => 
                           REGISTERS_9_26_port, QN => n17451);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n3889, CK => CLK, Q => 
                           REGISTERS_9_25_port, QN => n17212);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n3888, CK => CLK, Q => 
                           REGISTERS_9_24_port, QN => n17213);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n3887, CK => CLK, Q => 
                           REGISTERS_9_23_port, QN => n17452);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n3886, CK => CLK, Q => 
                           REGISTERS_9_22_port, QN => n17214);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n3885, CK => CLK, Q => 
                           REGISTERS_9_21_port, QN => n17453);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n3884, CK => CLK, Q => 
                           REGISTERS_9_20_port, QN => n17215);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n3883, CK => CLK, Q => 
                           REGISTERS_9_19_port, QN => n17454);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n3882, CK => CLK, Q => 
                           REGISTERS_9_18_port, QN => n17216);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n3881, CK => CLK, Q => 
                           REGISTERS_9_17_port, QN => n17217);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n3880, CK => CLK, Q => 
                           REGISTERS_9_16_port, QN => n17218);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n3879, CK => CLK, Q => 
                           REGISTERS_9_15_port, QN => n18491);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n3878, CK => CLK, Q => 
                           REGISTERS_9_14_port, QN => n18492);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n3877, CK => CLK, Q => 
                           REGISTERS_9_13_port, QN => n18133);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n3876, CK => CLK, Q => 
                           REGISTERS_9_12_port, QN => n18493);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n3875, CK => CLK, Q => 
                           REGISTERS_9_11_port, QN => n18134);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n3874, CK => CLK, Q => 
                           REGISTERS_9_10_port, QN => n18135);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n3873, CK => CLK, Q => 
                           REGISTERS_9_9_port, QN => n18136);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n3872, CK => CLK, Q => 
                           REGISTERS_9_8_port, QN => n18494);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n3871, CK => CLK, Q => 
                           REGISTERS_9_7_port, QN => n18137);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n3870, CK => CLK, Q => 
                           REGISTERS_9_6_port, QN => n18138);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n3869, CK => CLK, Q => 
                           REGISTERS_9_5_port, QN => n18495);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n3868, CK => CLK, Q => 
                           REGISTERS_9_4_port, QN => n18807);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n3867, CK => CLK, Q => 
                           REGISTERS_9_3_port, QN => n18139);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n3866, CK => CLK, Q => 
                           REGISTERS_9_2_port, QN => n18140);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n3865, CK => CLK, Q => 
                           REGISTERS_9_1_port, QN => n18141);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n3864, CK => CLK, Q => 
                           REGISTERS_9_0_port, QN => n18142);
   REGISTERS_reg_10_63_inst : DFF_X1 port map( D => n3863, CK => CLK, Q => 
                           REGISTERS_10_63_port, QN => n16888);
   REGISTERS_reg_10_62_inst : DFF_X1 port map( D => n3862, CK => CLK, Q => 
                           REGISTERS_10_62_port, QN => n18496);
   REGISTERS_reg_10_61_inst : DFF_X1 port map( D => n3861, CK => CLK, Q => 
                           REGISTERS_10_61_port, QN => n18143);
   REGISTERS_reg_10_60_inst : DFF_X1 port map( D => n3860, CK => CLK, Q => 
                           REGISTERS_10_60_port, QN => n18144);
   REGISTERS_reg_10_59_inst : DFF_X1 port map( D => n3859, CK => CLK, Q => 
                           REGISTERS_10_59_port, QN => n18145);
   REGISTERS_reg_10_58_inst : DFF_X1 port map( D => n3858, CK => n13730, Q => 
                           REGISTERS_10_58_port, QN => n18146);
   REGISTERS_reg_10_57_inst : DFF_X1 port map( D => n3857, CK => CLK, Q => 
                           REGISTERS_10_57_port, QN => n18147);
   REGISTERS_reg_10_56_inst : DFF_X1 port map( D => n3856, CK => n13730, Q => 
                           REGISTERS_10_56_port, QN => n18148);
   REGISTERS_reg_10_55_inst : DFF_X1 port map( D => n3855, CK => CLK, Q => 
                           REGISTERS_10_55_port, QN => n18497);
   REGISTERS_reg_10_54_inst : DFF_X1 port map( D => n3854, CK => CLK, Q => 
                           REGISTERS_10_54_port, QN => n18498);
   REGISTERS_reg_10_53_inst : DFF_X1 port map( D => n3853, CK => CLK, Q => 
                           REGISTERS_10_53_port, QN => n18149);
   REGISTERS_reg_10_52_inst : DFF_X1 port map( D => n3852, CK => CLK, Q => 
                           REGISTERS_10_52_port, QN => n18499);
   REGISTERS_reg_10_51_inst : DFF_X1 port map( D => n3851, CK => CLK, Q => 
                           REGISTERS_10_51_port, QN => n18150);
   REGISTERS_reg_10_50_inst : DFF_X1 port map( D => n3850, CK => CLK, Q => 
                           REGISTERS_10_50_port, QN => n18500);
   REGISTERS_reg_10_49_inst : DFF_X1 port map( D => n3849, CK => CLK, Q => 
                           REGISTERS_10_49_port, QN => n18151);
   REGISTERS_reg_10_48_inst : DFF_X1 port map( D => n3848, CK => CLK, Q => 
                           REGISTERS_10_48_port, QN => n18501);
   REGISTERS_reg_10_47_inst : DFF_X1 port map( D => n3847, CK => CLK, Q => 
                           REGISTERS_10_47_port, QN => n18502);
   REGISTERS_reg_10_46_inst : DFF_X1 port map( D => n3846, CK => CLK, Q => 
                           REGISTERS_10_46_port, QN => n18503);
   REGISTERS_reg_10_45_inst : DFF_X1 port map( D => n3845, CK => CLK, Q => 
                           REGISTERS_10_45_port, QN => n18504);
   REGISTERS_reg_10_44_inst : DFF_X1 port map( D => n3844, CK => CLK, Q => 
                           REGISTERS_10_44_port, QN => n18808);
   REGISTERS_reg_10_43_inst : DFF_X1 port map( D => n3843, CK => CLK, Q => 
                           REGISTERS_10_43_port, QN => n18505);
   REGISTERS_reg_10_42_inst : DFF_X1 port map( D => n3842, CK => CLK, Q => 
                           REGISTERS_10_42_port, QN => n18506);
   REGISTERS_reg_10_41_inst : DFF_X1 port map( D => n3841, CK => CLK, Q => 
                           REGISTERS_10_41_port, QN => n18809);
   REGISTERS_reg_10_40_inst : DFF_X1 port map( D => n3840, CK => CLK, Q => 
                           REGISTERS_10_40_port, QN => n18152);
   REGISTERS_reg_10_39_inst : DFF_X1 port map( D => n3839, CK => CLK, Q => 
                           REGISTERS_10_39_port, QN => n18507);
   REGISTERS_reg_10_38_inst : DFF_X1 port map( D => n3838, CK => CLK, Q => 
                           REGISTERS_10_38_port, QN => n18508);
   REGISTERS_reg_10_37_inst : DFF_X1 port map( D => n3837, CK => CLK, Q => 
                           REGISTERS_10_37_port, QN => n18509);
   REGISTERS_reg_10_36_inst : DFF_X1 port map( D => n3836, CK => CLK, Q => 
                           REGISTERS_10_36_port, QN => n18510);
   REGISTERS_reg_10_35_inst : DFF_X1 port map( D => n3835, CK => CLK, Q => 
                           REGISTERS_10_35_port, QN => n18153);
   REGISTERS_reg_10_34_inst : DFF_X1 port map( D => n3834, CK => CLK, Q => 
                           REGISTERS_10_34_port, QN => n18511);
   REGISTERS_reg_10_33_inst : DFF_X1 port map( D => n3833, CK => CLK, Q => 
                           REGISTERS_10_33_port, QN => n18512);
   REGISTERS_reg_10_32_inst : DFF_X1 port map( D => n3832, CK => CLK, Q => 
                           REGISTERS_10_32_port, QN => n18810);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n3831, CK => CLK, Q => 
                           REGISTERS_10_31_port, QN => n18154);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n3830, CK => CLK, Q => 
                           REGISTERS_10_30_port, QN => n18513);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n3829, CK => CLK, Q => 
                           REGISTERS_10_29_port, QN => n18155);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n3828, CK => CLK, Q => 
                           REGISTERS_10_28_port, QN => n18514);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n3827, CK => CLK, Q => 
                           REGISTERS_10_27_port, QN => n17219);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n3826, CK => CLK, Q => 
                           REGISTERS_10_26_port, QN => n17220);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n3825, CK => CLK, Q => 
                           REGISTERS_10_25_port, QN => n17824);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n3824, CK => CLK, Q => 
                           REGISTERS_10_24_port, QN => n17221);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n3823, CK => CLK, Q => 
                           REGISTERS_10_23_port, QN => n17455);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n3822, CK => CLK, Q => 
                           REGISTERS_10_22_port, QN => n17825);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n3821, CK => CLK, Q => 
                           REGISTERS_10_21_port, QN => n17826);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n3820, CK => CLK, Q => 
                           REGISTERS_10_20_port, QN => n17456);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n3819, CK => CLK, Q => 
                           REGISTERS_10_19_port, QN => n17457);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n3818, CK => CLK, Q => 
                           REGISTERS_10_18_port, QN => n17458);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n3817, CK => CLK, Q => 
                           REGISTERS_10_17_port, QN => n17459);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n3816, CK => CLK, Q => 
                           REGISTERS_10_16_port, QN => n17222);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n3815, CK => CLK, Q => 
                           REGISTERS_10_15_port, QN => n18156);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n3814, CK => CLK, Q => 
                           REGISTERS_10_14_port, QN => n18515);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n3813, CK => n13730, Q => 
                           REGISTERS_10_13_port, QN => n18516);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n3812, CK => CLK, Q => 
                           REGISTERS_10_12_port, QN => n18517);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n3811, CK => CLK, Q => 
                           REGISTERS_10_11_port, QN => n18811);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n3810, CK => CLK, Q => 
                           REGISTERS_10_10_port, QN => n18157);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n3809, CK => CLK, Q => 
                           REGISTERS_10_9_port, QN => n18158);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n3808, CK => n13730, Q => 
                           REGISTERS_10_8_port, QN => n18518);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n3807, CK => CLK, Q => 
                           REGISTERS_10_7_port, QN => n18519);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n3806, CK => CLK, Q => 
                           REGISTERS_10_6_port, QN => n18520);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n3805, CK => CLK, Q => 
                           REGISTERS_10_5_port, QN => n18812);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n3804, CK => CLK, Q => 
                           REGISTERS_10_4_port, QN => n18159);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n3803, CK => CLK, Q => 
                           REGISTERS_10_3_port, QN => n18160);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n3802, CK => CLK, Q => 
                           REGISTERS_10_2_port, QN => n18521);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n3801, CK => CLK, Q => 
                           REGISTERS_10_1_port, QN => n18161);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n3800, CK => CLK, Q => 
                           REGISTERS_10_0_port, QN => n18522);
   REGISTERS_reg_11_63_inst : DFF_X1 port map( D => n3799, CK => CLK, Q => 
                           REGISTERS_11_63_port, QN => n16965);
   REGISTERS_reg_11_62_inst : DFF_X1 port map( D => n3798, CK => CLK, Q => 
                           REGISTERS_11_62_port, QN => n18523);
   REGISTERS_reg_11_61_inst : DFF_X1 port map( D => n3797, CK => CLK, Q => 
                           REGISTERS_11_61_port, QN => n18813);
   REGISTERS_reg_11_60_inst : DFF_X1 port map( D => n3796, CK => CLK, Q => 
                           REGISTERS_11_60_port, QN => n18162);
   REGISTERS_reg_11_59_inst : DFF_X1 port map( D => n3795, CK => CLK, Q => 
                           REGISTERS_11_59_port, QN => n18814);
   REGISTERS_reg_11_58_inst : DFF_X1 port map( D => n3794, CK => CLK, Q => 
                           REGISTERS_11_58_port, QN => n18163);
   REGISTERS_reg_11_57_inst : DFF_X1 port map( D => n3793, CK => CLK, Q => 
                           REGISTERS_11_57_port, QN => n18524);
   REGISTERS_reg_11_56_inst : DFF_X1 port map( D => n3792, CK => CLK, Q => 
                           REGISTERS_11_56_port, QN => n18815);
   REGISTERS_reg_11_55_inst : DFF_X1 port map( D => n3791, CK => CLK, Q => 
                           REGISTERS_11_55_port, QN => n18816);
   REGISTERS_reg_11_54_inst : DFF_X1 port map( D => n3790, CK => CLK, Q => 
                           REGISTERS_11_54_port, QN => n18164);
   REGISTERS_reg_11_53_inst : DFF_X1 port map( D => n3789, CK => CLK, Q => 
                           REGISTERS_11_53_port, QN => n18525);
   REGISTERS_reg_11_52_inst : DFF_X1 port map( D => n3788, CK => CLK, Q => 
                           REGISTERS_11_52_port, QN => n18165);
   REGISTERS_reg_11_51_inst : DFF_X1 port map( D => n3787, CK => CLK, Q => 
                           REGISTERS_11_51_port, QN => n18526);
   REGISTERS_reg_11_50_inst : DFF_X1 port map( D => n3786, CK => CLK, Q => 
                           REGISTERS_11_50_port, QN => n18527);
   REGISTERS_reg_11_49_inst : DFF_X1 port map( D => n3785, CK => CLK, Q => 
                           REGISTERS_11_49_port, QN => n18166);
   REGISTERS_reg_11_48_inst : DFF_X1 port map( D => n3784, CK => CLK, Q => 
                           REGISTERS_11_48_port, QN => n18528);
   REGISTERS_reg_11_47_inst : DFF_X1 port map( D => n3783, CK => CLK, Q => 
                           REGISTERS_11_47_port, QN => n18529);
   REGISTERS_reg_11_46_inst : DFF_X1 port map( D => n3782, CK => CLK, Q => 
                           REGISTERS_11_46_port, QN => n18530);
   REGISTERS_reg_11_45_inst : DFF_X1 port map( D => n3781, CK => CLK, Q => 
                           REGISTERS_11_45_port, QN => n18531);
   REGISTERS_reg_11_44_inst : DFF_X1 port map( D => n3780, CK => n13730, Q => 
                           REGISTERS_11_44_port, QN => n18167);
   REGISTERS_reg_11_43_inst : DFF_X1 port map( D => n3779, CK => CLK, Q => 
                           REGISTERS_11_43_port, QN => n18817);
   REGISTERS_reg_11_42_inst : DFF_X1 port map( D => n3778, CK => CLK, Q => 
                           REGISTERS_11_42_port, QN => n18532);
   REGISTERS_reg_11_41_inst : DFF_X1 port map( D => n3777, CK => CLK, Q => 
                           REGISTERS_11_41_port, QN => n18818);
   REGISTERS_reg_11_40_inst : DFF_X1 port map( D => n3776, CK => CLK, Q => 
                           REGISTERS_11_40_port, QN => n18168);
   REGISTERS_reg_11_39_inst : DFF_X1 port map( D => n3775, CK => CLK, Q => 
                           REGISTERS_11_39_port, QN => n18533);
   REGISTERS_reg_11_38_inst : DFF_X1 port map( D => n3774, CK => CLK, Q => 
                           REGISTERS_11_38_port, QN => n18819);
   REGISTERS_reg_11_37_inst : DFF_X1 port map( D => n3773, CK => CLK, Q => 
                           REGISTERS_11_37_port, QN => n18534);
   REGISTERS_reg_11_36_inst : DFF_X1 port map( D => n3772, CK => CLK, Q => 
                           REGISTERS_11_36_port, QN => n18169);
   REGISTERS_reg_11_35_inst : DFF_X1 port map( D => n3771, CK => CLK, Q => 
                           REGISTERS_11_35_port, QN => n18535);
   REGISTERS_reg_11_34_inst : DFF_X1 port map( D => n3770, CK => CLK, Q => 
                           REGISTERS_11_34_port, QN => n18536);
   REGISTERS_reg_11_33_inst : DFF_X1 port map( D => n3769, CK => CLK, Q => 
                           REGISTERS_11_33_port, QN => n18820);
   REGISTERS_reg_11_32_inst : DFF_X1 port map( D => n3768, CK => CLK, Q => 
                           REGISTERS_11_32_port, QN => n18170);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n3767, CK => CLK, Q => 
                           REGISTERS_11_31_port, QN => n18821);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n3766, CK => CLK, Q => 
                           REGISTERS_11_30_port, QN => n18171);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n3765, CK => CLK, Q => 
                           REGISTERS_11_29_port, QN => n18822);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n3764, CK => CLK, Q => 
                           REGISTERS_11_28_port, QN => n18172);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n3763, CK => CLK, Q => 
                           REGISTERS_11_27_port, QN => n17223);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n3762, CK => CLK, Q => 
                           REGISTERS_11_26_port, QN => n17460);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n3761, CK => CLK, Q => 
                           REGISTERS_11_25_port, QN => n17461);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n3760, CK => CLK, Q => 
                           REGISTERS_11_24_port, QN => n17827);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n3759, CK => CLK, Q => 
                           REGISTERS_11_23_port, QN => n17828);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n3758, CK => CLK, Q => 
                           REGISTERS_11_22_port, QN => n17462);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n3757, CK => CLK, Q => 
                           REGISTERS_11_21_port, QN => n17829);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n3756, CK => CLK, Q => 
                           REGISTERS_11_20_port, QN => n17224);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n3755, CK => CLK, Q => 
                           REGISTERS_11_19_port, QN => n17463);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n3754, CK => CLK, Q => 
                           REGISTERS_11_18_port, QN => n17464);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n3753, CK => CLK, Q => 
                           REGISTERS_11_17_port, QN => n17225);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n3752, CK => CLK, Q => 
                           REGISTERS_11_16_port, QN => n17465);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n3751, CK => CLK, Q => 
                           REGISTERS_11_15_port, QN => n18173);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n3750, CK => CLK, Q => 
                           REGISTERS_11_14_port, QN => n18174);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n3749, CK => CLK, Q => 
                           REGISTERS_11_13_port, QN => n18537);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n3748, CK => CLK, Q => 
                           REGISTERS_11_12_port, QN => n18823);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n3747, CK => CLK, Q => 
                           REGISTERS_11_11_port, QN => n18538);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n3746, CK => CLK, Q => 
                           REGISTERS_11_10_port, QN => n18824);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n3745, CK => CLK, Q => 
                           REGISTERS_11_9_port, QN => n18825);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n3744, CK => CLK, Q => 
                           REGISTERS_11_8_port, QN => n18826);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n3743, CK => CLK, Q => 
                           REGISTERS_11_7_port, QN => n18827);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n3742, CK => CLK, Q => 
                           REGISTERS_11_6_port, QN => n18175);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n3741, CK => CLK, Q => 
                           REGISTERS_11_5_port, QN => n18828);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n3740, CK => CLK, Q => 
                           REGISTERS_11_4_port, QN => n18539);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n3739, CK => CLK, Q => 
                           REGISTERS_11_3_port, QN => n18540);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n3738, CK => CLK, Q => 
                           REGISTERS_11_2_port, QN => n18541);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n3737, CK => CLK, Q => 
                           REGISTERS_11_1_port, QN => n18829);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n3736, CK => CLK, Q => 
                           REGISTERS_11_0_port, QN => n18176);
   REGISTERS_reg_12_63_inst : DFF_X1 port map( D => n3735, CK => CLK, Q => 
                           REGISTERS_12_63_port, QN => n17226);
   REGISTERS_reg_12_62_inst : DFF_X1 port map( D => n3734, CK => CLK, Q => 
                           REGISTERS_12_62_port, QN => n17227);
   REGISTERS_reg_12_61_inst : DFF_X1 port map( D => n3733, CK => CLK, Q => 
                           REGISTERS_12_61_port, QN => n17228);
   REGISTERS_reg_12_60_inst : DFF_X1 port map( D => n3732, CK => CLK, Q => 
                           REGISTERS_12_60_port, QN => n17466);
   REGISTERS_reg_12_59_inst : DFF_X1 port map( D => n3731, CK => CLK, Q => 
                           REGISTERS_12_59_port, QN => n17467);
   REGISTERS_reg_12_58_inst : DFF_X1 port map( D => n3730, CK => CLK, Q => 
                           REGISTERS_12_58_port, QN => n17468);
   REGISTERS_reg_12_57_inst : DFF_X1 port map( D => n3729, CK => CLK, Q => 
                           REGISTERS_12_57_port, QN => n17469);
   REGISTERS_reg_12_56_inst : DFF_X1 port map( D => n3728, CK => CLK, Q => 
                           REGISTERS_12_56_port, QN => n17470);
   REGISTERS_reg_12_55_inst : DFF_X1 port map( D => n3727, CK => CLK, Q => 
                           REGISTERS_12_55_port, QN => n17471);
   REGISTERS_reg_12_54_inst : DFF_X1 port map( D => n3726, CK => CLK, Q => 
                           REGISTERS_12_54_port, QN => n17830);
   REGISTERS_reg_12_53_inst : DFF_X1 port map( D => n3725, CK => CLK, Q => 
                           REGISTERS_12_53_port, QN => n17472);
   REGISTERS_reg_12_52_inst : DFF_X1 port map( D => n3724, CK => CLK, Q => 
                           REGISTERS_12_52_port, QN => n17473);
   REGISTERS_reg_12_51_inst : DFF_X1 port map( D => n3723, CK => CLK, Q => 
                           REGISTERS_12_51_port, QN => n18542);
   REGISTERS_reg_12_50_inst : DFF_X1 port map( D => n3722, CK => CLK, Q => 
                           REGISTERS_12_50_port, QN => n18543);
   REGISTERS_reg_12_49_inst : DFF_X1 port map( D => n3721, CK => CLK, Q => 
                           REGISTERS_12_49_port, QN => n18177);
   REGISTERS_reg_12_48_inst : DFF_X1 port map( D => n3720, CK => CLK, Q => 
                           REGISTERS_12_48_port, QN => n18830);
   REGISTERS_reg_12_47_inst : DFF_X1 port map( D => n3719, CK => CLK, Q => 
                           REGISTERS_12_47_port, QN => n18178);
   REGISTERS_reg_12_46_inst : DFF_X1 port map( D => n3718, CK => CLK, Q => 
                           REGISTERS_12_46_port, QN => n18544);
   REGISTERS_reg_12_45_inst : DFF_X1 port map( D => n3717, CK => CLK, Q => 
                           REGISTERS_12_45_port, QN => n18831);
   REGISTERS_reg_12_44_inst : DFF_X1 port map( D => n3716, CK => CLK, Q => 
                           REGISTERS_12_44_port, QN => n18545);
   REGISTERS_reg_12_43_inst : DFF_X1 port map( D => n3715, CK => CLK, Q => 
                           REGISTERS_12_43_port, QN => n18546);
   REGISTERS_reg_12_42_inst : DFF_X1 port map( D => n3714, CK => CLK, Q => 
                           REGISTERS_12_42_port, QN => n18179);
   REGISTERS_reg_12_41_inst : DFF_X1 port map( D => n3713, CK => CLK, Q => 
                           REGISTERS_12_41_port, QN => n18547);
   REGISTERS_reg_12_40_inst : DFF_X1 port map( D => n3712, CK => CLK, Q => 
                           REGISTERS_12_40_port, QN => n18548);
   REGISTERS_reg_12_39_inst : DFF_X1 port map( D => n3711, CK => CLK, Q => 
                           REGISTERS_12_39_port, QN => n18549);
   REGISTERS_reg_12_38_inst : DFF_X1 port map( D => n3710, CK => CLK, Q => 
                           REGISTERS_12_38_port, QN => n18180);
   REGISTERS_reg_12_37_inst : DFF_X1 port map( D => n3709, CK => CLK, Q => 
                           REGISTERS_12_37_port, QN => n18550);
   REGISTERS_reg_12_36_inst : DFF_X1 port map( D => n3708, CK => CLK, Q => 
                           REGISTERS_12_36_port, QN => n18551);
   REGISTERS_reg_12_35_inst : DFF_X1 port map( D => n3707, CK => CLK, Q => 
                           REGISTERS_12_35_port, QN => n18552);
   REGISTERS_reg_12_34_inst : DFF_X1 port map( D => n3706, CK => CLK, Q => 
                           REGISTERS_12_34_port, QN => n18832);
   REGISTERS_reg_12_33_inst : DFF_X1 port map( D => n3705, CK => CLK, Q => 
                           REGISTERS_12_33_port, QN => n18833);
   REGISTERS_reg_12_32_inst : DFF_X1 port map( D => n3704, CK => CLK, Q => 
                           REGISTERS_12_32_port, QN => n18553);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n3703, CK => CLK, Q => 
                           REGISTERS_12_31_port, QN => n18554);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n3702, CK => CLK, Q => 
                           REGISTERS_12_30_port, QN => n18555);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n3701, CK => CLK, Q => 
                           REGISTERS_12_29_port, QN => n18834);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n3700, CK => CLK, Q => 
                           REGISTERS_12_28_port, QN => n18556);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n3699, CK => CLK, Q => 
                           REGISTERS_12_27_port, QN => n17831);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n3698, CK => CLK, Q => 
                           REGISTERS_12_26_port, QN => n17474);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n3697, CK => CLK, Q => 
                           REGISTERS_12_25_port, QN => n17475);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n3696, CK => CLK, Q => 
                           REGISTERS_12_24_port, QN => n17229);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n3695, CK => CLK, Q => 
                           REGISTERS_12_23_port, QN => n17832);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n3694, CK => CLK, Q => 
                           REGISTERS_12_22_port, QN => n17476);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n3693, CK => CLK, Q => 
                           REGISTERS_12_21_port, QN => n17477);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n3692, CK => CLK, Q => 
                           REGISTERS_12_20_port, QN => n17478);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n3691, CK => CLK, Q => 
                           REGISTERS_12_19_port, QN => n17230);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n3690, CK => CLK, Q => 
                           REGISTERS_12_18_port, QN => n17479);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n3689, CK => CLK, Q => 
                           REGISTERS_12_17_port, QN => n17833);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n3688, CK => CLK, Q => 
                           REGISTERS_12_16_port, QN => n17834);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n3687, CK => CLK, Q => 
                           REGISTERS_12_15_port, QN => n18557);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n3686, CK => CLK, Q => 
                           REGISTERS_12_14_port, QN => n18835);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n3685, CK => CLK, Q => 
                           REGISTERS_12_13_port, QN => n18558);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n3684, CK => n13730, Q => 
                           REGISTERS_12_12_port, QN => n18836);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n3683, CK => CLK, Q => 
                           REGISTERS_12_11_port, QN => n18559);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n3682, CK => CLK, Q => 
                           REGISTERS_12_10_port, QN => n18837);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n3681, CK => CLK, Q => 
                           REGISTERS_12_9_port, QN => n18560);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n3680, CK => CLK, Q => 
                           REGISTERS_12_8_port, QN => n18561);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n3679, CK => CLK, Q => 
                           REGISTERS_12_7_port, QN => n18562);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n3678, CK => CLK, Q => 
                           REGISTERS_12_6_port, QN => n18838);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n3677, CK => CLK, Q => 
                           REGISTERS_12_5_port, QN => n18181);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n3676, CK => CLK, Q => 
                           REGISTERS_12_4_port, QN => n18182);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n3675, CK => CLK, Q => 
                           REGISTERS_12_3_port, QN => n18183);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n3674, CK => CLK, Q => 
                           REGISTERS_12_2_port, QN => n18563);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n3673, CK => CLK, Q => 
                           REGISTERS_12_1_port, QN => n18184);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n3672, CK => CLK, Q => 
                           REGISTERS_12_0_port, QN => n18185);
   REGISTERS_reg_13_63_inst : DFF_X1 port map( D => n3671, CK => CLK, Q => 
                           REGISTERS_13_63_port, QN => n17231);
   REGISTERS_reg_13_62_inst : DFF_X1 port map( D => n3670, CK => n13730, Q => 
                           REGISTERS_13_62_port, QN => n17835);
   REGISTERS_reg_13_61_inst : DFF_X1 port map( D => n3669, CK => CLK, Q => 
                           REGISTERS_13_61_port, QN => n17836);
   REGISTERS_reg_13_60_inst : DFF_X1 port map( D => n3668, CK => CLK, Q => 
                           REGISTERS_13_60_port, QN => n17837);
   REGISTERS_reg_13_59_inst : DFF_X1 port map( D => n3667, CK => CLK, Q => 
                           REGISTERS_13_59_port, QN => n17838);
   REGISTERS_reg_13_58_inst : DFF_X1 port map( D => n3666, CK => CLK, Q => 
                           REGISTERS_13_58_port, QN => n17839);
   REGISTERS_reg_13_57_inst : DFF_X1 port map( D => n3665, CK => CLK, Q => 
                           REGISTERS_13_57_port, QN => n17480);
   REGISTERS_reg_13_56_inst : DFF_X1 port map( D => n3664, CK => CLK, Q => 
                           REGISTERS_13_56_port, QN => n17840);
   REGISTERS_reg_13_55_inst : DFF_X1 port map( D => n3663, CK => CLK, Q => 
                           REGISTERS_13_55_port, QN => n17481);
   REGISTERS_reg_13_54_inst : DFF_X1 port map( D => n3662, CK => CLK, Q => 
                           REGISTERS_13_54_port, QN => n17482);
   REGISTERS_reg_13_53_inst : DFF_X1 port map( D => n3661, CK => CLK, Q => 
                           REGISTERS_13_53_port, QN => n17841);
   REGISTERS_reg_13_52_inst : DFF_X1 port map( D => n3660, CK => CLK, Q => 
                           REGISTERS_13_52_port, QN => n17842);
   REGISTERS_reg_13_51_inst : DFF_X1 port map( D => n3659, CK => CLK, Q => 
                           REGISTERS_13_51_port, QN => n18564);
   REGISTERS_reg_13_50_inst : DFF_X1 port map( D => n3658, CK => CLK, Q => 
                           REGISTERS_13_50_port, QN => n18839);
   REGISTERS_reg_13_49_inst : DFF_X1 port map( D => n3657, CK => CLK, Q => 
                           REGISTERS_13_49_port, QN => n18840);
   REGISTERS_reg_13_48_inst : DFF_X1 port map( D => n3656, CK => CLK, Q => 
                           REGISTERS_13_48_port, QN => n18841);
   REGISTERS_reg_13_47_inst : DFF_X1 port map( D => n3655, CK => CLK, Q => 
                           REGISTERS_13_47_port, QN => n18842);
   REGISTERS_reg_13_46_inst : DFF_X1 port map( D => n3654, CK => CLK, Q => 
                           REGISTERS_13_46_port, QN => n18843);
   REGISTERS_reg_13_45_inst : DFF_X1 port map( D => n3653, CK => CLK, Q => 
                           REGISTERS_13_45_port, QN => n18844);
   REGISTERS_reg_13_44_inst : DFF_X1 port map( D => n3652, CK => CLK, Q => 
                           REGISTERS_13_44_port, QN => n18565);
   REGISTERS_reg_13_43_inst : DFF_X1 port map( D => n3651, CK => CLK, Q => 
                           REGISTERS_13_43_port, QN => n18566);
   REGISTERS_reg_13_42_inst : DFF_X1 port map( D => n3650, CK => CLK, Q => 
                           REGISTERS_13_42_port, QN => n18845);
   REGISTERS_reg_13_41_inst : DFF_X1 port map( D => n3649, CK => CLK, Q => 
                           REGISTERS_13_41_port, QN => n18567);
   REGISTERS_reg_13_40_inst : DFF_X1 port map( D => n3648, CK => CLK, Q => 
                           REGISTERS_13_40_port, QN => n18846);
   REGISTERS_reg_13_39_inst : DFF_X1 port map( D => n3647, CK => CLK, Q => 
                           REGISTERS_13_39_port, QN => n18568);
   REGISTERS_reg_13_38_inst : DFF_X1 port map( D => n3646, CK => CLK, Q => 
                           REGISTERS_13_38_port, QN => n18847);
   REGISTERS_reg_13_37_inst : DFF_X1 port map( D => n3645, CK => CLK, Q => 
                           REGISTERS_13_37_port, QN => n18569);
   REGISTERS_reg_13_36_inst : DFF_X1 port map( D => n3644, CK => CLK, Q => 
                           REGISTERS_13_36_port, QN => n18570);
   REGISTERS_reg_13_35_inst : DFF_X1 port map( D => n3643, CK => CLK, Q => 
                           REGISTERS_13_35_port, QN => n18848);
   REGISTERS_reg_13_34_inst : DFF_X1 port map( D => n3642, CK => CLK, Q => 
                           REGISTERS_13_34_port, QN => n18849);
   REGISTERS_reg_13_33_inst : DFF_X1 port map( D => n3641, CK => CLK, Q => 
                           REGISTERS_13_33_port, QN => n18571);
   REGISTERS_reg_13_32_inst : DFF_X1 port map( D => n3640, CK => CLK, Q => 
                           REGISTERS_13_32_port, QN => n18850);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n3639, CK => CLK, Q => 
                           REGISTERS_13_31_port, QN => n18572);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n3638, CK => CLK, Q => 
                           REGISTERS_13_30_port, QN => n18851);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n3637, CK => CLK, Q => 
                           REGISTERS_13_29_port, QN => n18573);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n3636, CK => CLK, Q => 
                           REGISTERS_13_28_port, QN => n18574);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n3635, CK => CLK, Q => 
                           REGISTERS_13_27_port, QN => n17232);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n3634, CK => CLK, Q => 
                           REGISTERS_13_26_port, QN => n17843);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n3633, CK => CLK, Q => 
                           REGISTERS_13_25_port, QN => n17233);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n3632, CK => CLK, Q => 
                           REGISTERS_13_24_port, QN => n17483);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n3631, CK => CLK, Q => 
                           REGISTERS_13_23_port, QN => n17484);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n3630, CK => CLK, Q => 
                           REGISTERS_13_22_port, QN => n17844);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n3629, CK => CLK, Q => 
                           REGISTERS_13_21_port, QN => n17485);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n3628, CK => CLK, Q => 
                           REGISTERS_13_20_port, QN => n17845);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n3627, CK => CLK, Q => 
                           REGISTERS_13_19_port, QN => n17846);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n3626, CK => CLK, Q => 
                           REGISTERS_13_18_port, QN => n17847);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n3625, CK => CLK, Q => 
                           REGISTERS_13_17_port, QN => n17486);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n3624, CK => CLK, Q => 
                           REGISTERS_13_16_port, QN => n17487);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n3623, CK => CLK, Q => 
                           REGISTERS_13_15_port, QN => n18575);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n3622, CK => CLK, Q => 
                           REGISTERS_13_14_port, QN => n18576);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n3621, CK => CLK, Q => 
                           REGISTERS_13_13_port, QN => n18577);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n3620, CK => CLK, Q => 
                           REGISTERS_13_12_port, QN => n18578);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n3619, CK => CLK, Q => 
                           REGISTERS_13_11_port, QN => n18579);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n3618, CK => CLK, Q => 
                           REGISTERS_13_10_port, QN => n18580);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n3617, CK => CLK, Q => 
                           REGISTERS_13_9_port, QN => n18852);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n3616, CK => CLK, Q => 
                           REGISTERS_13_8_port, QN => n18581);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n3615, CK => CLK, Q => 
                           REGISTERS_13_7_port, QN => n18853);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n3614, CK => CLK, Q => 
                           REGISTERS_13_6_port, QN => n18582);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n3613, CK => CLK, Q => 
                           REGISTERS_13_5_port, QN => n18854);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n3612, CK => CLK, Q => 
                           REGISTERS_13_4_port, QN => n18855);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n3611, CK => CLK, Q => 
                           REGISTERS_13_3_port, QN => n18856);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n3610, CK => CLK, Q => 
                           REGISTERS_13_2_port, QN => n18857);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n3609, CK => CLK, Q => 
                           REGISTERS_13_1_port, QN => n18858);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n3608, CK => CLK, Q => 
                           REGISTERS_13_0_port, QN => n18859);
   REGISTERS_reg_14_63_inst : DFF_X1 port map( D => n3607, CK => CLK, Q => 
                           REGISTERS_14_63_port, QN => n17171);
   REGISTERS_reg_14_62_inst : DFF_X1 port map( D => n3606, CK => CLK, Q => 
                           REGISTERS_14_62_port, QN => n17234);
   REGISTERS_reg_14_61_inst : DFF_X1 port map( D => n3605, CK => CLK, Q => 
                           REGISTERS_14_61_port, QN => n17488);
   REGISTERS_reg_14_60_inst : DFF_X1 port map( D => n3604, CK => CLK, Q => 
                           REGISTERS_14_60_port, QN => n17489);
   REGISTERS_reg_14_59_inst : DFF_X1 port map( D => n3603, CK => CLK, Q => 
                           REGISTERS_14_59_port, QN => n17490);
   REGISTERS_reg_14_58_inst : DFF_X1 port map( D => n3602, CK => CLK, Q => 
                           REGISTERS_14_58_port, QN => n17491);
   REGISTERS_reg_14_57_inst : DFF_X1 port map( D => n3601, CK => CLK, Q => 
                           REGISTERS_14_57_port, QN => n17235);
   REGISTERS_reg_14_56_inst : DFF_X1 port map( D => n3600, CK => CLK, Q => 
                           REGISTERS_14_56_port, QN => n17236);
   REGISTERS_reg_14_55_inst : DFF_X1 port map( D => n3599, CK => CLK, Q => 
                           REGISTERS_14_55_port, QN => n17237);
   REGISTERS_reg_14_54_inst : DFF_X1 port map( D => n3598, CK => CLK, Q => 
                           REGISTERS_14_54_port, QN => n17238);
   REGISTERS_reg_14_53_inst : DFF_X1 port map( D => n3597, CK => CLK, Q => 
                           REGISTERS_14_53_port, QN => n17492);
   REGISTERS_reg_14_52_inst : DFF_X1 port map( D => n3596, CK => CLK, Q => 
                           REGISTERS_14_52_port, QN => n17493);
   REGISTERS_reg_14_51_inst : DFF_X1 port map( D => n3595, CK => CLK, Q => 
                           REGISTERS_14_51_port, QN => n18583);
   REGISTERS_reg_14_50_inst : DFF_X1 port map( D => n3594, CK => CLK, Q => 
                           REGISTERS_14_50_port, QN => n18584);
   REGISTERS_reg_14_49_inst : DFF_X1 port map( D => n3593, CK => CLK, Q => 
                           REGISTERS_14_49_port, QN => n18585);
   REGISTERS_reg_14_48_inst : DFF_X1 port map( D => n3592, CK => CLK, Q => 
                           REGISTERS_14_48_port, QN => n18586);
   REGISTERS_reg_14_47_inst : DFF_X1 port map( D => n3591, CK => CLK, Q => 
                           REGISTERS_14_47_port, QN => n18587);
   REGISTERS_reg_14_46_inst : DFF_X1 port map( D => n3590, CK => CLK, Q => 
                           REGISTERS_14_46_port, QN => n18186);
   REGISTERS_reg_14_45_inst : DFF_X1 port map( D => n3589, CK => CLK, Q => 
                           REGISTERS_14_45_port, QN => n18187);
   REGISTERS_reg_14_44_inst : DFF_X1 port map( D => n3588, CK => CLK, Q => 
                           REGISTERS_14_44_port, QN => n18188);
   REGISTERS_reg_14_43_inst : DFF_X1 port map( D => n3587, CK => CLK, Q => 
                           REGISTERS_14_43_port, QN => n18588);
   REGISTERS_reg_14_42_inst : DFF_X1 port map( D => n3586, CK => CLK, Q => 
                           REGISTERS_14_42_port, QN => n18189);
   REGISTERS_reg_14_41_inst : DFF_X1 port map( D => n3585, CK => CLK, Q => 
                           REGISTERS_14_41_port, QN => n18860);
   REGISTERS_reg_14_40_inst : DFF_X1 port map( D => n3584, CK => CLK, Q => 
                           REGISTERS_14_40_port, QN => n18589);
   REGISTERS_reg_14_39_inst : DFF_X1 port map( D => n3583, CK => CLK, Q => 
                           REGISTERS_14_39_port, QN => n18190);
   REGISTERS_reg_14_38_inst : DFF_X1 port map( D => n3582, CK => CLK, Q => 
                           REGISTERS_14_38_port, QN => n18191);
   REGISTERS_reg_14_37_inst : DFF_X1 port map( D => n3581, CK => CLK, Q => 
                           REGISTERS_14_37_port, QN => n18192);
   REGISTERS_reg_14_36_inst : DFF_X1 port map( D => n3580, CK => CLK, Q => 
                           REGISTERS_14_36_port, QN => n18193);
   REGISTERS_reg_14_35_inst : DFF_X1 port map( D => n3579, CK => CLK, Q => 
                           REGISTERS_14_35_port, QN => n18590);
   REGISTERS_reg_14_34_inst : DFF_X1 port map( D => n3578, CK => CLK, Q => 
                           REGISTERS_14_34_port, QN => n18591);
   REGISTERS_reg_14_33_inst : DFF_X1 port map( D => n3577, CK => CLK, Q => 
                           REGISTERS_14_33_port, QN => n18592);
   REGISTERS_reg_14_32_inst : DFF_X1 port map( D => n3576, CK => CLK, Q => 
                           REGISTERS_14_32_port, QN => n18194);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n3575, CK => CLK, Q => 
                           REGISTERS_14_31_port, QN => n18593);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n3574, CK => CLK, Q => 
                           REGISTERS_14_30_port, QN => n18195);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n3573, CK => CLK, Q => 
                           REGISTERS_14_29_port, QN => n18594);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n3572, CK => CLK, Q => 
                           REGISTERS_14_28_port, QN => n18595);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n3571, CK => CLK, Q => 
                           REGISTERS_14_27_port, QN => n17494);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n3570, CK => CLK, Q => 
                           REGISTERS_14_26_port, QN => n17495);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n3569, CK => CLK, Q => 
                           REGISTERS_14_25_port, QN => n17496);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n3568, CK => CLK, Q => 
                           REGISTERS_14_24_port, QN => n17848);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n3567, CK => CLK, Q => 
                           REGISTERS_14_23_port, QN => n17497);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n3566, CK => CLK, Q => 
                           REGISTERS_14_22_port, QN => n17498);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n3565, CK => CLK, Q => 
                           REGISTERS_14_21_port, QN => n17239);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n3564, CK => CLK, Q => 
                           REGISTERS_14_20_port, QN => n17499);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n3563, CK => CLK, Q => 
                           REGISTERS_14_19_port, QN => n17500);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n3562, CK => CLK, Q => 
                           REGISTERS_14_18_port, QN => n17240);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n3561, CK => CLK, Q => 
                           REGISTERS_14_17_port, QN => n17241);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n3560, CK => CLK, Q => 
                           REGISTERS_14_16_port, QN => n17849);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n3559, CK => CLK, Q => 
                           REGISTERS_14_15_port, QN => n18596);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n3558, CK => CLK, Q => 
                           REGISTERS_14_14_port, QN => n18597);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n3557, CK => CLK, Q => 
                           REGISTERS_14_13_port, QN => n18196);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n3556, CK => CLK, Q => 
                           REGISTERS_14_12_port, QN => n18598);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n3555, CK => CLK, Q => 
                           REGISTERS_14_11_port, QN => n18599);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n3554, CK => CLK, Q => 
                           REGISTERS_14_10_port, QN => n18600);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n3553, CK => CLK, Q => 
                           REGISTERS_14_9_port, QN => n18197);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n3552, CK => CLK, Q => 
                           REGISTERS_14_8_port, QN => n18198);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n3551, CK => CLK, Q => 
                           REGISTERS_14_7_port, QN => n18199);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n3550, CK => CLK, Q => 
                           REGISTERS_14_6_port, QN => n18601);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n3549, CK => CLK, Q => 
                           REGISTERS_14_5_port, QN => n18200);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n3548, CK => CLK, Q => 
                           REGISTERS_14_4_port, QN => n18602);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n3547, CK => CLK, Q => 
                           REGISTERS_14_3_port, QN => n18603);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n3546, CK => CLK, Q => 
                           REGISTERS_14_2_port, QN => n18604);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n3545, CK => CLK, Q => 
                           REGISTERS_14_1_port, QN => n18201);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n3544, CK => CLK, Q => 
                           REGISTERS_14_0_port, QN => n18202);
   REGISTERS_reg_15_63_inst : DFF_X1 port map( D => n3543, CK => CLK, Q => 
                           REGISTERS_15_63_port, QN => n17501);
   REGISTERS_reg_15_62_inst : DFF_X1 port map( D => n3542, CK => CLK, Q => 
                           REGISTERS_15_62_port, QN => n17850);
   REGISTERS_reg_15_61_inst : DFF_X1 port map( D => n3541, CK => CLK, Q => 
                           REGISTERS_15_61_port, QN => n17502);
   REGISTERS_reg_15_60_inst : DFF_X1 port map( D => n3540, CK => CLK, Q => 
                           REGISTERS_15_60_port, QN => n17851);
   REGISTERS_reg_15_59_inst : DFF_X1 port map( D => n3539, CK => CLK, Q => 
                           REGISTERS_15_59_port, QN => n17503);
   REGISTERS_reg_15_58_inst : DFF_X1 port map( D => n3538, CK => CLK, Q => 
                           REGISTERS_15_58_port, QN => n17504);
   REGISTERS_reg_15_57_inst : DFF_X1 port map( D => n3537, CK => CLK, Q => 
                           REGISTERS_15_57_port, QN => n17242);
   REGISTERS_reg_15_56_inst : DFF_X1 port map( D => n3536, CK => CLK, Q => 
                           REGISTERS_15_56_port, QN => n17243);
   REGISTERS_reg_15_55_inst : DFF_X1 port map( D => n3535, CK => CLK, Q => 
                           REGISTERS_15_55_port, QN => n17852);
   REGISTERS_reg_15_54_inst : DFF_X1 port map( D => n3534, CK => CLK, Q => 
                           REGISTERS_15_54_port, QN => n17244);
   REGISTERS_reg_15_53_inst : DFF_X1 port map( D => n3533, CK => CLK, Q => 
                           REGISTERS_15_53_port, QN => n17505);
   REGISTERS_reg_15_52_inst : DFF_X1 port map( D => n3532, CK => CLK, Q => 
                           REGISTERS_15_52_port, QN => n17853);
   REGISTERS_reg_15_51_inst : DFF_X1 port map( D => n3531, CK => CLK, Q => 
                           REGISTERS_15_51_port, QN => n18605);
   REGISTERS_reg_15_50_inst : DFF_X1 port map( D => n3530, CK => CLK, Q => 
                           REGISTERS_15_50_port, QN => n18203);
   REGISTERS_reg_15_49_inst : DFF_X1 port map( D => n3529, CK => CLK, Q => 
                           REGISTERS_15_49_port, QN => n18606);
   REGISTERS_reg_15_48_inst : DFF_X1 port map( D => n3528, CK => CLK, Q => 
                           REGISTERS_15_48_port, QN => n18607);
   REGISTERS_reg_15_47_inst : DFF_X1 port map( D => n3527, CK => CLK, Q => 
                           REGISTERS_15_47_port, QN => n18608);
   REGISTERS_reg_15_46_inst : DFF_X1 port map( D => n3526, CK => n13730, Q => 
                           REGISTERS_15_46_port, QN => n18861);
   REGISTERS_reg_15_45_inst : DFF_X1 port map( D => n3525, CK => CLK, Q => 
                           REGISTERS_15_45_port, QN => n18204);
   REGISTERS_reg_15_44_inst : DFF_X1 port map( D => n3524, CK => CLK, Q => 
                           REGISTERS_15_44_port, QN => n18205);
   REGISTERS_reg_15_43_inst : DFF_X1 port map( D => n3523, CK => CLK, Q => 
                           REGISTERS_15_43_port, QN => n18862);
   REGISTERS_reg_15_42_inst : DFF_X1 port map( D => n3522, CK => CLK, Q => 
                           REGISTERS_15_42_port, QN => n18609);
   REGISTERS_reg_15_41_inst : DFF_X1 port map( D => n3521, CK => CLK, Q => 
                           REGISTERS_15_41_port, QN => n18610);
   REGISTERS_reg_15_40_inst : DFF_X1 port map( D => n3520, CK => CLK, Q => 
                           REGISTERS_15_40_port, QN => n18863);
   REGISTERS_reg_15_39_inst : DFF_X1 port map( D => n3519, CK => CLK, Q => 
                           REGISTERS_15_39_port, QN => n18864);
   REGISTERS_reg_15_38_inst : DFF_X1 port map( D => n3518, CK => CLK, Q => 
                           REGISTERS_15_38_port, QN => n18206);
   REGISTERS_reg_15_37_inst : DFF_X1 port map( D => n3517, CK => CLK, Q => 
                           REGISTERS_15_37_port, QN => n18611);
   REGISTERS_reg_15_36_inst : DFF_X1 port map( D => n3516, CK => CLK, Q => 
                           REGISTERS_15_36_port, QN => n18207);
   REGISTERS_reg_15_35_inst : DFF_X1 port map( D => n3515, CK => CLK, Q => 
                           REGISTERS_15_35_port, QN => n18208);
   REGISTERS_reg_15_34_inst : DFF_X1 port map( D => n3514, CK => CLK, Q => 
                           REGISTERS_15_34_port, QN => n18612);
   REGISTERS_reg_15_33_inst : DFF_X1 port map( D => n3513, CK => CLK, Q => 
                           REGISTERS_15_33_port, QN => n18865);
   REGISTERS_reg_15_32_inst : DFF_X1 port map( D => n3512, CK => CLK, Q => 
                           REGISTERS_15_32_port, QN => n18866);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n3511, CK => CLK, Q => 
                           REGISTERS_15_31_port, QN => n18613);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n3510, CK => CLK, Q => 
                           REGISTERS_15_30_port, QN => n18614);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n3509, CK => CLK, Q => 
                           REGISTERS_15_29_port, QN => n18615);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n3508, CK => CLK, Q => 
                           REGISTERS_15_28_port, QN => n18867);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n3507, CK => CLK, Q => 
                           REGISTERS_15_27_port, QN => n17506);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n3506, CK => CLK, Q => 
                           REGISTERS_15_26_port, QN => n17507);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n3505, CK => CLK, Q => 
                           REGISTERS_15_25_port, QN => n17245);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n3504, CK => CLK, Q => 
                           REGISTERS_15_24_port, QN => n17508);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n3503, CK => CLK, Q => 
                           REGISTERS_15_23_port, QN => n17509);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n3502, CK => CLK, Q => 
                           REGISTERS_15_22_port, QN => n17854);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n3501, CK => CLK, Q => 
                           REGISTERS_15_21_port, QN => n17510);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n3500, CK => CLK, Q => 
                           REGISTERS_15_20_port, QN => n17246);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n3499, CK => CLK, Q => 
                           REGISTERS_15_19_port, QN => n17855);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n3498, CK => CLK, Q => 
                           REGISTERS_15_18_port, QN => n17511);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n3497, CK => CLK, Q => 
                           REGISTERS_15_17_port, QN => n17512);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n3496, CK => CLK, Q => 
                           REGISTERS_15_16_port, QN => n17856);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n3495, CK => CLK, Q => 
                           REGISTERS_15_15_port, QN => n18616);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n3494, CK => CLK, Q => 
                           REGISTERS_15_14_port, QN => n18209);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n3493, CK => CLK, Q => 
                           REGISTERS_15_13_port, QN => n18868);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n3492, CK => CLK, Q => 
                           REGISTERS_15_12_port, QN => n18617);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n3491, CK => CLK, Q => 
                           REGISTERS_15_11_port, QN => n18210);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n3490, CK => CLK, Q => 
                           REGISTERS_15_10_port, QN => n18211);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n3489, CK => CLK, Q => 
                           REGISTERS_15_9_port, QN => n18212);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n3488, CK => CLK, Q => 
                           REGISTERS_15_8_port, QN => n18618);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n3487, CK => CLK, Q => 
                           REGISTERS_15_7_port, QN => n18213);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n3486, CK => CLK, Q => 
                           REGISTERS_15_6_port, QN => n18869);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n3485, CK => CLK, Q => 
                           REGISTERS_15_5_port, QN => n18619);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n3484, CK => CLK, Q => 
                           REGISTERS_15_4_port, QN => n18870);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n3483, CK => CLK, Q => 
                           REGISTERS_15_3_port, QN => n18620);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n3482, CK => CLK, Q => 
                           REGISTERS_15_2_port, QN => n18871);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n3481, CK => CLK, Q => 
                           REGISTERS_15_1_port, QN => n18621);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n3480, CK => CLK, Q => 
                           REGISTERS_15_0_port, QN => n18622);
   REGISTERS_reg_16_63_inst : DFF_X1 port map( D => n3479, CK => CLK, Q => 
                           REGISTERS_16_63_port, QN => n17513);
   REGISTERS_reg_16_62_inst : DFF_X1 port map( D => n3478, CK => CLK, Q => 
                           REGISTERS_16_62_port, QN => n17514);
   REGISTERS_reg_16_61_inst : DFF_X1 port map( D => n3477, CK => CLK, Q => 
                           REGISTERS_16_61_port, QN => n17515);
   REGISTERS_reg_16_60_inst : DFF_X1 port map( D => n3476, CK => CLK, Q => 
                           REGISTERS_16_60_port, QN => n17247);
   REGISTERS_reg_16_59_inst : DFF_X1 port map( D => n3475, CK => CLK, Q => 
                           REGISTERS_16_59_port, QN => n17248);
   REGISTERS_reg_16_58_inst : DFF_X1 port map( D => n3474, CK => CLK, Q => 
                           REGISTERS_16_58_port, QN => n17516);
   REGISTERS_reg_16_57_inst : DFF_X1 port map( D => n3473, CK => CLK, Q => 
                           REGISTERS_16_57_port, QN => n17517);
   REGISTERS_reg_16_56_inst : DFF_X1 port map( D => n3472, CK => n13730, Q => 
                           REGISTERS_16_56_port, QN => n17857);
   REGISTERS_reg_16_55_inst : DFF_X1 port map( D => n3471, CK => CLK, Q => 
                           REGISTERS_16_55_port, QN => n17518);
   REGISTERS_reg_16_54_inst : DFF_X1 port map( D => n3470, CK => CLK, Q => 
                           REGISTERS_16_54_port, QN => n17858);
   REGISTERS_reg_16_53_inst : DFF_X1 port map( D => n3469, CK => CLK, Q => 
                           REGISTERS_16_53_port, QN => n17519);
   REGISTERS_reg_16_52_inst : DFF_X1 port map( D => n3468, CK => CLK, Q => 
                           REGISTERS_16_52_port, QN => n17520);
   REGISTERS_reg_16_51_inst : DFF_X1 port map( D => n3467, CK => CLK, Q => 
                           REGISTERS_16_51_port, QN => n18214);
   REGISTERS_reg_16_50_inst : DFF_X1 port map( D => n3466, CK => CLK, Q => 
                           REGISTERS_16_50_port, QN => n18215);
   REGISTERS_reg_16_49_inst : DFF_X1 port map( D => n3465, CK => CLK, Q => 
                           REGISTERS_16_49_port, QN => n18623);
   REGISTERS_reg_16_48_inst : DFF_X1 port map( D => n3464, CK => CLK, Q => 
                           REGISTERS_16_48_port, QN => n18216);
   REGISTERS_reg_16_47_inst : DFF_X1 port map( D => n3463, CK => CLK, Q => 
                           REGISTERS_16_47_port, QN => n18624);
   REGISTERS_reg_16_46_inst : DFF_X1 port map( D => n3462, CK => CLK, Q => 
                           REGISTERS_16_46_port, QN => n18625);
   REGISTERS_reg_16_45_inst : DFF_X1 port map( D => n3461, CK => CLK, Q => 
                           REGISTERS_16_45_port, QN => n18872);
   REGISTERS_reg_16_44_inst : DFF_X1 port map( D => n3460, CK => CLK, Q => 
                           REGISTERS_16_44_port, QN => n18217);
   REGISTERS_reg_16_43_inst : DFF_X1 port map( D => n3459, CK => CLK, Q => 
                           REGISTERS_16_43_port, QN => n18626);
   REGISTERS_reg_16_42_inst : DFF_X1 port map( D => n3458, CK => CLK, Q => 
                           REGISTERS_16_42_port, QN => n18627);
   REGISTERS_reg_16_41_inst : DFF_X1 port map( D => n3457, CK => CLK, Q => 
                           REGISTERS_16_41_port, QN => n18628);
   REGISTERS_reg_16_40_inst : DFF_X1 port map( D => n3456, CK => CLK, Q => 
                           REGISTERS_16_40_port, QN => n18218);
   REGISTERS_reg_16_39_inst : DFF_X1 port map( D => n3455, CK => CLK, Q => 
                           REGISTERS_16_39_port, QN => n18219);
   REGISTERS_reg_16_38_inst : DFF_X1 port map( D => n3454, CK => CLK, Q => 
                           REGISTERS_16_38_port, QN => n18629);
   REGISTERS_reg_16_37_inst : DFF_X1 port map( D => n3453, CK => CLK, Q => 
                           REGISTERS_16_37_port, QN => n18873);
   REGISTERS_reg_16_36_inst : DFF_X1 port map( D => n3452, CK => CLK, Q => 
                           REGISTERS_16_36_port, QN => n18630);
   REGISTERS_reg_16_35_inst : DFF_X1 port map( D => n3451, CK => CLK, Q => 
                           REGISTERS_16_35_port, QN => n18220);
   REGISTERS_reg_16_34_inst : DFF_X1 port map( D => n3450, CK => CLK, Q => 
                           REGISTERS_16_34_port, QN => n18221);
   REGISTERS_reg_16_33_inst : DFF_X1 port map( D => n3449, CK => CLK, Q => 
                           REGISTERS_16_33_port, QN => n18631);
   REGISTERS_reg_16_32_inst : DFF_X1 port map( D => n3448, CK => CLK, Q => 
                           REGISTERS_16_32_port, QN => n18632);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n3447, CK => CLK, Q => 
                           REGISTERS_16_31_port, QN => n18874);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n3446, CK => CLK, Q => 
                           REGISTERS_16_30_port, QN => n18633);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n3445, CK => CLK, Q => 
                           REGISTERS_16_29_port, QN => n18222);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n3444, CK => CLK, Q => 
                           REGISTERS_16_28_port, QN => n18634);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n3443, CK => CLK, Q => 
                           REGISTERS_16_27_port, QN => n17249);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n3442, CK => CLK, Q => 
                           REGISTERS_16_26_port, QN => n17859);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n3441, CK => CLK, Q => 
                           REGISTERS_16_25_port, QN => n17521);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n3440, CK => CLK, Q => 
                           REGISTERS_16_24_port, QN => n17522);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n3439, CK => CLK, Q => 
                           REGISTERS_16_23_port, QN => n17860);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n3438, CK => CLK, Q => 
                           REGISTERS_16_22_port, QN => n17861);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n3437, CK => CLK, Q => 
                           REGISTERS_16_21_port, QN => n17523);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n3436, CK => CLK, Q => 
                           REGISTERS_16_20_port, QN => n17524);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n3435, CK => CLK, Q => 
                           REGISTERS_16_19_port, QN => n17525);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n3434, CK => CLK, Q => 
                           REGISTERS_16_18_port, QN => n17526);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n3433, CK => CLK, Q => 
                           REGISTERS_16_17_port, QN => n17527);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n3432, CK => CLK, Q => 
                           REGISTERS_16_16_port, QN => n17250);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n3431, CK => CLK, Q => 
                           REGISTERS_16_15_port, QN => n18223);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n3430, CK => CLK, Q => 
                           REGISTERS_16_14_port, QN => n18635);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n3429, CK => CLK, Q => 
                           REGISTERS_16_13_port, QN => n18224);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n3428, CK => CLK, Q => 
                           REGISTERS_16_12_port, QN => n18225);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n3427, CK => CLK, Q => 
                           REGISTERS_16_11_port, QN => n18636);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n3426, CK => CLK, Q => 
                           REGISTERS_16_10_port, QN => n18637);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n3425, CK => CLK, Q => 
                           REGISTERS_16_9_port, QN => n18875);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n3424, CK => CLK, Q => 
                           REGISTERS_16_8_port, QN => n18876);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n3423, CK => CLK, Q => 
                           REGISTERS_16_7_port, QN => n18226);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n3422, CK => CLK, Q => 
                           REGISTERS_16_6_port, QN => n18227);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n3421, CK => CLK, Q => 
                           REGISTERS_16_5_port, QN => n18228);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n3420, CK => CLK, Q => 
                           REGISTERS_16_4_port, QN => n18638);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n3419, CK => CLK, Q => 
                           REGISTERS_16_3_port, QN => n18639);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n3418, CK => CLK, Q => 
                           REGISTERS_16_2_port, QN => n18640);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n3417, CK => CLK, Q => 
                           REGISTERS_16_1_port, QN => n18641);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n3416, CK => CLK, Q => 
                           REGISTERS_16_0_port, QN => n18229);
   REGISTERS_reg_17_63_inst : DFF_X1 port map( D => n3415, CK => CLK, Q => 
                           REGISTERS_17_63_port, QN => n17251);
   REGISTERS_reg_17_62_inst : DFF_X1 port map( D => n3414, CK => CLK, Q => 
                           REGISTERS_17_62_port, QN => n17862);
   REGISTERS_reg_17_61_inst : DFF_X1 port map( D => n3413, CK => CLK, Q => 
                           REGISTERS_17_61_port, QN => n17528);
   REGISTERS_reg_17_60_inst : DFF_X1 port map( D => n3412, CK => CLK, Q => 
                           REGISTERS_17_60_port, QN => n17529);
   REGISTERS_reg_17_59_inst : DFF_X1 port map( D => n3411, CK => CLK, Q => 
                           REGISTERS_17_59_port, QN => n17530);
   REGISTERS_reg_17_58_inst : DFF_X1 port map( D => n3410, CK => CLK, Q => 
                           REGISTERS_17_58_port, QN => n17531);
   REGISTERS_reg_17_57_inst : DFF_X1 port map( D => n3409, CK => CLK, Q => 
                           REGISTERS_17_57_port, QN => n17863);
   REGISTERS_reg_17_56_inst : DFF_X1 port map( D => n3408, CK => CLK, Q => 
                           REGISTERS_17_56_port, QN => n17864);
   REGISTERS_reg_17_55_inst : DFF_X1 port map( D => n3407, CK => CLK, Q => 
                           REGISTERS_17_55_port, QN => n17532);
   REGISTERS_reg_17_54_inst : DFF_X1 port map( D => n3406, CK => CLK, Q => 
                           REGISTERS_17_54_port, QN => n17865);
   REGISTERS_reg_17_53_inst : DFF_X1 port map( D => n3405, CK => CLK, Q => 
                           REGISTERS_17_53_port, QN => n17533);
   REGISTERS_reg_17_52_inst : DFF_X1 port map( D => n3404, CK => CLK, Q => 
                           REGISTERS_17_52_port, QN => n17866);
   REGISTERS_reg_17_51_inst : DFF_X1 port map( D => n3403, CK => CLK, Q => 
                           REGISTERS_17_51_port, QN => n18877);
   REGISTERS_reg_17_50_inst : DFF_X1 port map( D => n3402, CK => CLK, Q => 
                           REGISTERS_17_50_port, QN => n18878);
   REGISTERS_reg_17_49_inst : DFF_X1 port map( D => n3401, CK => CLK, Q => 
                           REGISTERS_17_49_port, QN => n18879);
   REGISTERS_reg_17_48_inst : DFF_X1 port map( D => n3400, CK => CLK, Q => 
                           REGISTERS_17_48_port, QN => n18880);
   REGISTERS_reg_17_47_inst : DFF_X1 port map( D => n3399, CK => CLK, Q => 
                           REGISTERS_17_47_port, QN => n18881);
   REGISTERS_reg_17_46_inst : DFF_X1 port map( D => n3398, CK => CLK, Q => 
                           REGISTERS_17_46_port, QN => n18882);
   REGISTERS_reg_17_45_inst : DFF_X1 port map( D => n3397, CK => CLK, Q => 
                           REGISTERS_17_45_port, QN => n18883);
   REGISTERS_reg_17_44_inst : DFF_X1 port map( D => n3396, CK => CLK, Q => 
                           REGISTERS_17_44_port, QN => n18884);
   REGISTERS_reg_17_43_inst : DFF_X1 port map( D => n3395, CK => CLK, Q => 
                           REGISTERS_17_43_port, QN => n18885);
   REGISTERS_reg_17_42_inst : DFF_X1 port map( D => n3394, CK => CLK, Q => 
                           REGISTERS_17_42_port, QN => n18642);
   REGISTERS_reg_17_41_inst : DFF_X1 port map( D => n3393, CK => CLK, Q => 
                           REGISTERS_17_41_port, QN => n18643);
   REGISTERS_reg_17_40_inst : DFF_X1 port map( D => n3392, CK => CLK, Q => 
                           REGISTERS_17_40_port, QN => n18644);
   REGISTERS_reg_17_39_inst : DFF_X1 port map( D => n3391, CK => CLK, Q => 
                           REGISTERS_17_39_port, QN => n18645);
   REGISTERS_reg_17_38_inst : DFF_X1 port map( D => n3390, CK => CLK, Q => 
                           REGISTERS_17_38_port, QN => n18646);
   REGISTERS_reg_17_37_inst : DFF_X1 port map( D => n3389, CK => CLK, Q => 
                           REGISTERS_17_37_port, QN => n18886);
   REGISTERS_reg_17_36_inst : DFF_X1 port map( D => n3388, CK => CLK, Q => 
                           REGISTERS_17_36_port, QN => n18647);
   REGISTERS_reg_17_35_inst : DFF_X1 port map( D => n3387, CK => CLK, Q => 
                           REGISTERS_17_35_port, QN => n18648);
   REGISTERS_reg_17_34_inst : DFF_X1 port map( D => n3386, CK => CLK, Q => 
                           REGISTERS_17_34_port, QN => n18649);
   REGISTERS_reg_17_33_inst : DFF_X1 port map( D => n3385, CK => CLK, Q => 
                           REGISTERS_17_33_port, QN => n18650);
   REGISTERS_reg_17_32_inst : DFF_X1 port map( D => n3384, CK => CLK, Q => 
                           REGISTERS_17_32_port, QN => n18887);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n3383, CK => CLK, Q => 
                           REGISTERS_17_31_port, QN => n18651);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n3382, CK => CLK, Q => 
                           REGISTERS_17_30_port, QN => n18888);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n3381, CK => CLK, Q => 
                           REGISTERS_17_29_port, QN => n18889);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n3380, CK => CLK, Q => 
                           REGISTERS_17_28_port, QN => n18890);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n3379, CK => CLK, Q => 
                           REGISTERS_17_27_port, QN => n17534);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n3378, CK => n13730, Q => 
                           REGISTERS_17_26_port, QN => n17252);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n3377, CK => CLK, Q => 
                           REGISTERS_17_25_port, QN => n17535);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n3376, CK => CLK, Q => 
                           REGISTERS_17_24_port, QN => n17253);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n3375, CK => CLK, Q => 
                           REGISTERS_17_23_port, QN => n17867);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n3374, CK => CLK, Q => 
                           REGISTERS_17_22_port, QN => n17536);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n3373, CK => CLK, Q => 
                           REGISTERS_17_21_port, QN => n17537);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n3372, CK => CLK, Q => 
                           REGISTERS_17_20_port, QN => n17538);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n3371, CK => CLK, Q => 
                           REGISTERS_17_19_port, QN => n17868);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n3370, CK => CLK, Q => 
                           REGISTERS_17_18_port, QN => n17539);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n3369, CK => CLK, Q => 
                           REGISTERS_17_17_port, QN => n17869);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n3368, CK => CLK, Q => 
                           REGISTERS_17_16_port, QN => n17540);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n3367, CK => CLK, Q => 
                           REGISTERS_17_15_port, QN => n18652);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n3366, CK => CLK, Q => 
                           REGISTERS_17_14_port, QN => n18653);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n3365, CK => CLK, Q => 
                           REGISTERS_17_13_port, QN => n18891);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n3364, CK => CLK, Q => 
                           REGISTERS_17_12_port, QN => n18654);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n3363, CK => CLK, Q => 
                           REGISTERS_17_11_port, QN => n18892);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n3362, CK => CLK, Q => 
                           REGISTERS_17_10_port, QN => n18893);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n3361, CK => CLK, Q => 
                           REGISTERS_17_9_port, QN => n18655);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n3360, CK => CLK, Q => 
                           REGISTERS_17_8_port, QN => n18656);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n3359, CK => CLK, Q => 
                           REGISTERS_17_7_port, QN => n18894);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n3358, CK => CLK, Q => 
                           REGISTERS_17_6_port, QN => n18895);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n3357, CK => CLK, Q => 
                           REGISTERS_17_5_port, QN => n18230);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n3356, CK => CLK, Q => 
                           REGISTERS_17_4_port, QN => n18896);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n3355, CK => CLK, Q => 
                           REGISTERS_17_3_port, QN => n18657);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n3354, CK => CLK, Q => 
                           REGISTERS_17_2_port, QN => n18658);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n3353, CK => CLK, Q => 
                           REGISTERS_17_1_port, QN => n18659);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n3352, CK => CLK, Q => 
                           REGISTERS_17_0_port, QN => n18897);
   REGISTERS_reg_18_63_inst : DFF_X1 port map( D => n3351, CK => CLK, Q => 
                           REGISTERS_18_63_port, QN => n17541);
   REGISTERS_reg_18_62_inst : DFF_X1 port map( D => n3350, CK => CLK, Q => 
                           REGISTERS_18_62_port, QN => n17870);
   REGISTERS_reg_18_61_inst : DFF_X1 port map( D => n3349, CK => CLK, Q => 
                           REGISTERS_18_61_port, QN => n17542);
   REGISTERS_reg_18_60_inst : DFF_X1 port map( D => n3348, CK => CLK, Q => 
                           REGISTERS_18_60_port, QN => n17543);
   REGISTERS_reg_18_59_inst : DFF_X1 port map( D => n3347, CK => CLK, Q => 
                           REGISTERS_18_59_port, QN => n17254);
   REGISTERS_reg_18_58_inst : DFF_X1 port map( D => n3346, CK => CLK, Q => 
                           REGISTERS_18_58_port, QN => n17544);
   REGISTERS_reg_18_57_inst : DFF_X1 port map( D => n3345, CK => CLK, Q => 
                           REGISTERS_18_57_port, QN => n17871);
   REGISTERS_reg_18_56_inst : DFF_X1 port map( D => n3344, CK => CLK, Q => 
                           REGISTERS_18_56_port, QN => n17255);
   REGISTERS_reg_18_55_inst : DFF_X1 port map( D => n3343, CK => CLK, Q => 
                           REGISTERS_18_55_port, QN => n17545);
   REGISTERS_reg_18_54_inst : DFF_X1 port map( D => n3342, CK => CLK, Q => 
                           REGISTERS_18_54_port, QN => n17872);
   REGISTERS_reg_18_53_inst : DFF_X1 port map( D => n3341, CK => CLK, Q => 
                           REGISTERS_18_53_port, QN => n17546);
   REGISTERS_reg_18_52_inst : DFF_X1 port map( D => n3340, CK => CLK, Q => 
                           REGISTERS_18_52_port, QN => n17873);
   REGISTERS_reg_18_51_inst : DFF_X1 port map( D => n3339, CK => CLK, Q => 
                           REGISTERS_18_51_port, QN => n18898);
   REGISTERS_reg_18_50_inst : DFF_X1 port map( D => n3338, CK => CLK, Q => 
                           REGISTERS_18_50_port, QN => n18660);
   REGISTERS_reg_18_49_inst : DFF_X1 port map( D => n3337, CK => CLK, Q => 
                           REGISTERS_18_49_port, QN => n18661);
   REGISTERS_reg_18_48_inst : DFF_X1 port map( D => n3336, CK => CLK, Q => 
                           REGISTERS_18_48_port, QN => n18231);
   REGISTERS_reg_18_47_inst : DFF_X1 port map( D => n3335, CK => CLK, Q => 
                           REGISTERS_18_47_port, QN => n18662);
   REGISTERS_reg_18_46_inst : DFF_X1 port map( D => n3334, CK => CLK, Q => 
                           REGISTERS_18_46_port, QN => n18899);
   REGISTERS_reg_18_45_inst : DFF_X1 port map( D => n3333, CK => CLK, Q => 
                           REGISTERS_18_45_port, QN => n18900);
   REGISTERS_reg_18_44_inst : DFF_X1 port map( D => n3332, CK => CLK, Q => 
                           REGISTERS_18_44_port, QN => n18901);
   REGISTERS_reg_18_43_inst : DFF_X1 port map( D => n3331, CK => CLK, Q => 
                           REGISTERS_18_43_port, QN => n18902);
   REGISTERS_reg_18_42_inst : DFF_X1 port map( D => n3330, CK => CLK, Q => 
                           REGISTERS_18_42_port, QN => n18663);
   REGISTERS_reg_18_41_inst : DFF_X1 port map( D => n3329, CK => CLK, Q => 
                           REGISTERS_18_41_port, QN => n18903);
   REGISTERS_reg_18_40_inst : DFF_X1 port map( D => n3328, CK => CLK, Q => 
                           REGISTERS_18_40_port, QN => n18664);
   REGISTERS_reg_18_39_inst : DFF_X1 port map( D => n3327, CK => CLK, Q => 
                           REGISTERS_18_39_port, QN => n18904);
   REGISTERS_reg_18_38_inst : DFF_X1 port map( D => n3326, CK => n13730, Q => 
                           REGISTERS_18_38_port, QN => n18905);
   REGISTERS_reg_18_37_inst : DFF_X1 port map( D => n3325, CK => CLK, Q => 
                           REGISTERS_18_37_port, QN => n18665);
   REGISTERS_reg_18_36_inst : DFF_X1 port map( D => n3324, CK => CLK, Q => 
                           REGISTERS_18_36_port, QN => n18906);
   REGISTERS_reg_18_35_inst : DFF_X1 port map( D => n3323, CK => CLK, Q => 
                           REGISTERS_18_35_port, QN => n18666);
   REGISTERS_reg_18_34_inst : DFF_X1 port map( D => n3322, CK => CLK, Q => 
                           REGISTERS_18_34_port, QN => n18667);
   REGISTERS_reg_18_33_inst : DFF_X1 port map( D => n3321, CK => CLK, Q => 
                           REGISTERS_18_33_port, QN => n18232);
   REGISTERS_reg_18_32_inst : DFF_X1 port map( D => n3320, CK => CLK, Q => 
                           REGISTERS_18_32_port, QN => n18907);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n3319, CK => CLK, Q => 
                           REGISTERS_18_31_port, QN => n18668);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n3318, CK => CLK, Q => 
                           REGISTERS_18_30_port, QN => n18908);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n3317, CK => CLK, Q => 
                           REGISTERS_18_29_port, QN => n18909);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n3316, CK => CLK, Q => 
                           REGISTERS_18_28_port, QN => n18910);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n3315, CK => CLK, Q => 
                           REGISTERS_18_27_port, QN => n17547);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n3314, CK => CLK, Q => 
                           REGISTERS_18_26_port, QN => n17548);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n3313, CK => CLK, Q => 
                           REGISTERS_18_25_port, QN => n17874);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n3312, CK => CLK, Q => 
                           REGISTERS_18_24_port, QN => n17875);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n3311, CK => CLK, Q => 
                           REGISTERS_18_23_port, QN => n17549);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n3310, CK => CLK, Q => 
                           REGISTERS_18_22_port, QN => n17550);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n3309, CK => CLK, Q => 
                           REGISTERS_18_21_port, QN => n17551);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n3308, CK => CLK, Q => 
                           REGISTERS_18_20_port, QN => n17876);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n3307, CK => CLK, Q => 
                           REGISTERS_18_19_port, QN => n17552);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n3306, CK => CLK, Q => 
                           REGISTERS_18_18_port, QN => n17553);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n3305, CK => CLK, Q => 
                           REGISTERS_18_17_port, QN => n17554);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n3304, CK => CLK, Q => 
                           REGISTERS_18_16_port, QN => n17877);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n3303, CK => CLK, Q => 
                           REGISTERS_18_15_port, QN => n18669);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n3302, CK => CLK, Q => 
                           REGISTERS_18_14_port, QN => n18670);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n3301, CK => CLK, Q => 
                           REGISTERS_18_13_port, QN => n18911);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n3300, CK => CLK, Q => 
                           REGISTERS_18_12_port, QN => n18671);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n3299, CK => CLK, Q => 
                           REGISTERS_18_11_port, QN => n18912);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n3298, CK => CLK, Q => 
                           REGISTERS_18_10_port, QN => n18672);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n3297, CK => CLK, Q => 
                           REGISTERS_18_9_port, QN => n18913);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n3296, CK => CLK, Q => 
                           REGISTERS_18_8_port, QN => n18673);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n3295, CK => CLK, Q => 
                           REGISTERS_18_7_port, QN => n18674);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n3294, CK => CLK, Q => 
                           REGISTERS_18_6_port, QN => n18675);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n3293, CK => CLK, Q => 
                           REGISTERS_18_5_port, QN => n18676);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n3292, CK => CLK, Q => 
                           REGISTERS_18_4_port, QN => n18677);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n3291, CK => CLK, Q => 
                           REGISTERS_18_3_port, QN => n18914);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n3290, CK => CLK, Q => 
                           REGISTERS_18_2_port, QN => n18915);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n3289, CK => n13730, Q => 
                           REGISTERS_18_1_port, QN => n18678);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n3288, CK => CLK, Q => 
                           REGISTERS_18_0_port, QN => n18916);
   REGISTERS_reg_19_63_inst : DFF_X1 port map( D => n3287, CK => CLK, Q => 
                           REGISTERS_19_63_port, QN => n17555);
   REGISTERS_reg_19_62_inst : DFF_X1 port map( D => n3286, CK => CLK, Q => 
                           REGISTERS_19_62_port, QN => n17556);
   REGISTERS_reg_19_61_inst : DFF_X1 port map( D => n3285, CK => CLK, Q => 
                           REGISTERS_19_61_port, QN => n17878);
   REGISTERS_reg_19_60_inst : DFF_X1 port map( D => n3284, CK => CLK, Q => 
                           REGISTERS_19_60_port, QN => n17557);
   REGISTERS_reg_19_59_inst : DFF_X1 port map( D => n3283, CK => CLK, Q => 
                           REGISTERS_19_59_port, QN => n17558);
   REGISTERS_reg_19_58_inst : DFF_X1 port map( D => n3282, CK => CLK, Q => 
                           REGISTERS_19_58_port, QN => n17879);
   REGISTERS_reg_19_57_inst : DFF_X1 port map( D => n3281, CK => CLK, Q => 
                           REGISTERS_19_57_port, QN => n17880);
   REGISTERS_reg_19_56_inst : DFF_X1 port map( D => n3280, CK => CLK, Q => 
                           REGISTERS_19_56_port, QN => n17881);
   REGISTERS_reg_19_55_inst : DFF_X1 port map( D => n3279, CK => CLK, Q => 
                           REGISTERS_19_55_port, QN => n17559);
   REGISTERS_reg_19_54_inst : DFF_X1 port map( D => n3278, CK => CLK, Q => 
                           REGISTERS_19_54_port, QN => n17882);
   REGISTERS_reg_19_53_inst : DFF_X1 port map( D => n3277, CK => CLK, Q => 
                           REGISTERS_19_53_port, QN => n17560);
   REGISTERS_reg_19_52_inst : DFF_X1 port map( D => n3276, CK => CLK, Q => 
                           REGISTERS_19_52_port, QN => n17561);
   REGISTERS_reg_19_51_inst : DFF_X1 port map( D => n3275, CK => CLK, Q => 
                           REGISTERS_19_51_port, QN => n18917);
   REGISTERS_reg_19_50_inst : DFF_X1 port map( D => n3274, CK => CLK, Q => 
                           REGISTERS_19_50_port, QN => n18679);
   REGISTERS_reg_19_49_inst : DFF_X1 port map( D => n3273, CK => CLK, Q => 
                           REGISTERS_19_49_port, QN => n18233);
   REGISTERS_reg_19_48_inst : DFF_X1 port map( D => n3272, CK => CLK, Q => 
                           REGISTERS_19_48_port, QN => n18680);
   REGISTERS_reg_19_47_inst : DFF_X1 port map( D => n3271, CK => CLK, Q => 
                           REGISTERS_19_47_port, QN => n18918);
   REGISTERS_reg_19_46_inst : DFF_X1 port map( D => n3270, CK => CLK, Q => 
                           REGISTERS_19_46_port, QN => n18681);
   REGISTERS_reg_19_45_inst : DFF_X1 port map( D => n3269, CK => CLK, Q => 
                           REGISTERS_19_45_port, QN => n18682);
   REGISTERS_reg_19_44_inst : DFF_X1 port map( D => n3268, CK => CLK, Q => 
                           REGISTERS_19_44_port, QN => n18683);
   REGISTERS_reg_19_43_inst : DFF_X1 port map( D => n3267, CK => CLK, Q => 
                           REGISTERS_19_43_port, QN => n18919);
   REGISTERS_reg_19_42_inst : DFF_X1 port map( D => n3266, CK => CLK, Q => 
                           REGISTERS_19_42_port, QN => n18920);
   REGISTERS_reg_19_41_inst : DFF_X1 port map( D => n3265, CK => CLK, Q => 
                           REGISTERS_19_41_port, QN => n18234);
   REGISTERS_reg_19_40_inst : DFF_X1 port map( D => n3264, CK => CLK, Q => 
                           REGISTERS_19_40_port, QN => n18235);
   REGISTERS_reg_19_39_inst : DFF_X1 port map( D => n3263, CK => CLK, Q => 
                           REGISTERS_19_39_port, QN => n18921);
   REGISTERS_reg_19_38_inst : DFF_X1 port map( D => n3262, CK => CLK, Q => 
                           REGISTERS_19_38_port, QN => n18684);
   REGISTERS_reg_19_37_inst : DFF_X1 port map( D => n3261, CK => CLK, Q => 
                           REGISTERS_19_37_port, QN => n18922);
   REGISTERS_reg_19_36_inst : DFF_X1 port map( D => n3260, CK => CLK, Q => 
                           REGISTERS_19_36_port, QN => n18923);
   REGISTERS_reg_19_35_inst : DFF_X1 port map( D => n3259, CK => CLK, Q => 
                           REGISTERS_19_35_port, QN => n18236);
   REGISTERS_reg_19_34_inst : DFF_X1 port map( D => n3258, CK => CLK, Q => 
                           REGISTERS_19_34_port, QN => n18685);
   REGISTERS_reg_19_33_inst : DFF_X1 port map( D => n3257, CK => CLK, Q => 
                           REGISTERS_19_33_port, QN => n18686);
   REGISTERS_reg_19_32_inst : DFF_X1 port map( D => n3256, CK => CLK, Q => 
                           REGISTERS_19_32_port, QN => n18687);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n3255, CK => CLK, Q => 
                           REGISTERS_19_31_port, QN => n18924);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n3254, CK => CLK, Q => 
                           REGISTERS_19_30_port, QN => n18237);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n3253, CK => CLK, Q => 
                           REGISTERS_19_29_port, QN => n18688);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n3252, CK => CLK, Q => 
                           REGISTERS_19_28_port, QN => n18689);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n3251, CK => CLK, Q => 
                           REGISTERS_19_27_port, QN => n17883);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n3250, CK => CLK, Q => 
                           REGISTERS_19_26_port, QN => n17562);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n3249, CK => CLK, Q => 
                           REGISTERS_19_25_port, QN => n17884);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n3248, CK => CLK, Q => 
                           REGISTERS_19_24_port, QN => n17563);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n3247, CK => CLK, Q => 
                           REGISTERS_19_23_port, QN => n17564);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n3246, CK => CLK, Q => 
                           REGISTERS_19_22_port, QN => n17256);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n3245, CK => CLK, Q => 
                           REGISTERS_19_21_port, QN => n17885);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n3244, CK => CLK, Q => 
                           REGISTERS_19_20_port, QN => n17565);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n3243, CK => CLK, Q => 
                           REGISTERS_19_19_port, QN => n17566);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n3242, CK => CLK, Q => 
                           REGISTERS_19_18_port, QN => n17567);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n3241, CK => CLK, Q => 
                           REGISTERS_19_17_port, QN => n17257);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n3240, CK => CLK, Q => 
                           REGISTERS_19_16_port, QN => n17568);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n3239, CK => CLK, Q => 
                           REGISTERS_19_15_port, QN => n18690);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n3238, CK => CLK, Q => 
                           REGISTERS_19_14_port, QN => n18925);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n3237, CK => CLK, Q => 
                           REGISTERS_19_13_port, QN => n18926);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n3236, CK => CLK, Q => 
                           REGISTERS_19_12_port, QN => n18238);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n3235, CK => CLK, Q => 
                           REGISTERS_19_11_port, QN => n18927);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n3234, CK => CLK, Q => 
                           REGISTERS_19_10_port, QN => n18691);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n3233, CK => CLK, Q => 
                           REGISTERS_19_9_port, QN => n18692);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n3232, CK => CLK, Q => 
                           REGISTERS_19_8_port, QN => n18693);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n3231, CK => CLK, Q => 
                           REGISTERS_19_7_port, QN => n18694);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n3230, CK => CLK, Q => 
                           REGISTERS_19_6_port, QN => n18239);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n3229, CK => CLK, Q => 
                           REGISTERS_19_5_port, QN => n18928);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n3228, CK => CLK, Q => 
                           REGISTERS_19_4_port, QN => n18695);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n3227, CK => CLK, Q => 
                           REGISTERS_19_3_port, QN => n18929);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n3226, CK => CLK, Q => 
                           REGISTERS_19_2_port, QN => n18696);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n3225, CK => CLK, Q => 
                           REGISTERS_19_1_port, QN => n18930);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n3224, CK => CLK, Q => 
                           REGISTERS_19_0_port, QN => n18697);
   REGISTERS_reg_20_63_inst : DFF_X1 port map( D => n3223, CK => CLK, Q => 
                           REGISTERS_20_63_port, QN => n18011);
   REGISTERS_reg_20_62_inst : DFF_X1 port map( D => n3222, CK => CLK, Q => 
                           REGISTERS_20_62_port, QN => n16966);
   REGISTERS_reg_20_61_inst : DFF_X1 port map( D => n3221, CK => CLK, Q => 
                           REGISTERS_20_61_port, QN => n16889);
   REGISTERS_reg_20_60_inst : DFF_X1 port map( D => n3220, CK => CLK, Q => 
                           REGISTERS_20_60_port, QN => n16967);
   REGISTERS_reg_20_59_inst : DFF_X1 port map( D => n3219, CK => CLK, Q => 
                           REGISTERS_20_59_port, QN => n16968);
   REGISTERS_reg_20_58_inst : DFF_X1 port map( D => n3218, CK => CLK, Q => 
                           REGISTERS_20_58_port, QN => n16969);
   REGISTERS_reg_20_57_inst : DFF_X1 port map( D => n3217, CK => CLK, Q => 
                           REGISTERS_20_57_port, QN => n17108);
   REGISTERS_reg_20_56_inst : DFF_X1 port map( D => n3216, CK => CLK, Q => 
                           REGISTERS_20_56_port, QN => n16970);
   REGISTERS_reg_20_55_inst : DFF_X1 port map( D => n3215, CK => CLK, Q => 
                           REGISTERS_20_55_port, QN => n16890);
   REGISTERS_reg_20_54_inst : DFF_X1 port map( D => n3214, CK => CLK, Q => 
                           REGISTERS_20_54_port, QN => n16891);
   REGISTERS_reg_20_53_inst : DFF_X1 port map( D => n3213, CK => CLK, Q => 
                           REGISTERS_20_53_port, QN => n17109);
   REGISTERS_reg_20_52_inst : DFF_X1 port map( D => n3212, CK => CLK, Q => 
                           REGISTERS_20_52_port, QN => n16892);
   REGISTERS_reg_20_51_inst : DFF_X1 port map( D => n3211, CK => CLK, Q => 
                           REGISTERS_20_51_port, QN => n17569);
   REGISTERS_reg_20_50_inst : DFF_X1 port map( D => n3210, CK => CLK, Q => 
                           REGISTERS_20_50_port, QN => n17570);
   REGISTERS_reg_20_49_inst : DFF_X1 port map( D => n3209, CK => CLK, Q => 
                           REGISTERS_20_49_port, QN => n17571);
   REGISTERS_reg_20_48_inst : DFF_X1 port map( D => n3208, CK => n13730, Q => 
                           REGISTERS_20_48_port, QN => n17572);
   REGISTERS_reg_20_47_inst : DFF_X1 port map( D => n3207, CK => CLK, Q => 
                           REGISTERS_20_47_port, QN => n17886);
   REGISTERS_reg_20_46_inst : DFF_X1 port map( D => n3206, CK => CLK, Q => 
                           REGISTERS_20_46_port, QN => n17258);
   REGISTERS_reg_20_45_inst : DFF_X1 port map( D => n3205, CK => CLK, Q => 
                           REGISTERS_20_45_port, QN => n17259);
   REGISTERS_reg_20_44_inst : DFF_X1 port map( D => n3204, CK => CLK, Q => 
                           REGISTERS_20_44_port, QN => n17887);
   REGISTERS_reg_20_43_inst : DFF_X1 port map( D => n3203, CK => CLK, Q => 
                           REGISTERS_20_43_port, QN => n17573);
   REGISTERS_reg_20_42_inst : DFF_X1 port map( D => n3202, CK => CLK, Q => 
                           REGISTERS_20_42_port, QN => n17574);
   REGISTERS_reg_20_41_inst : DFF_X1 port map( D => n3201, CK => CLK, Q => 
                           REGISTERS_20_41_port, QN => n17260);
   REGISTERS_reg_20_40_inst : DFF_X1 port map( D => n3200, CK => CLK, Q => 
                           REGISTERS_20_40_port, QN => n17888);
   REGISTERS_reg_20_39_inst : DFF_X1 port map( D => n3199, CK => CLK, Q => 
                           REGISTERS_20_39_port, QN => n17575);
   REGISTERS_reg_20_38_inst : DFF_X1 port map( D => n3198, CK => CLK, Q => 
                           REGISTERS_20_38_port, QN => n17261);
   REGISTERS_reg_20_37_inst : DFF_X1 port map( D => n3197, CK => CLK, Q => 
                           REGISTERS_20_37_port, QN => n17889);
   REGISTERS_reg_20_36_inst : DFF_X1 port map( D => n3196, CK => CLK, Q => 
                           REGISTERS_20_36_port, QN => n17262);
   REGISTERS_reg_20_35_inst : DFF_X1 port map( D => n3195, CK => CLK, Q => 
                           REGISTERS_20_35_port, QN => n17576);
   REGISTERS_reg_20_34_inst : DFF_X1 port map( D => n3194, CK => CLK, Q => 
                           REGISTERS_20_34_port, QN => n17263);
   REGISTERS_reg_20_33_inst : DFF_X1 port map( D => n3193, CK => n13730, Q => 
                           REGISTERS_20_33_port, QN => n17890);
   REGISTERS_reg_20_32_inst : DFF_X1 port map( D => n3192, CK => CLK, Q => 
                           REGISTERS_20_32_port, QN => n17577);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n3191, CK => CLK, Q => 
                           REGISTERS_20_31_port, QN => n17891);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n3190, CK => CLK, Q => 
                           REGISTERS_20_30_port, QN => n17892);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n3189, CK => CLK, Q => 
                           REGISTERS_20_29_port, QN => n17578);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n3188, CK => CLK, Q => 
                           REGISTERS_20_28_port, QN => n17579);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n3187, CK => CLK, Q => 
                           REGISTERS_20_27_port, QN => n16893);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n3186, CK => CLK, Q => 
                           REGISTERS_20_26_port, QN => n16971);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n3185, CK => CLK, Q => 
                           REGISTERS_20_25_port, QN => n16972);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n3184, CK => CLK, Q => 
                           REGISTERS_20_24_port, QN => n16973);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n3183, CK => CLK, Q => 
                           REGISTERS_20_23_port, QN => n16974);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n3182, CK => CLK, Q => 
                           REGISTERS_20_22_port, QN => n16894);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n3181, CK => CLK, Q => 
                           REGISTERS_20_21_port, QN => n16975);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n3180, CK => CLK, Q => 
                           REGISTERS_20_20_port, QN => n16976);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n3179, CK => CLK, Q => 
                           REGISTERS_20_19_port, QN => n16977);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n3178, CK => CLK, Q => 
                           REGISTERS_20_18_port, QN => n17110);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n3177, CK => n13730, Q => 
                           REGISTERS_20_17_port, QN => n17111);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n3176, CK => CLK, Q => 
                           REGISTERS_20_16_port, QN => n16978);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n3175, CK => CLK, Q => 
                           REGISTERS_20_15_port, QN => n17893);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n3174, CK => CLK, Q => 
                           REGISTERS_20_14_port, QN => n17894);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n3173, CK => CLK, Q => 
                           REGISTERS_20_13_port, QN => n17580);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n3172, CK => CLK, Q => 
                           REGISTERS_20_12_port, QN => n17581);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n3171, CK => CLK, Q => 
                           REGISTERS_20_11_port, QN => n17895);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n3170, CK => CLK, Q => 
                           REGISTERS_20_10_port, QN => n17264);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n3169, CK => CLK, Q => 
                           REGISTERS_20_9_port, QN => n17582);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n3168, CK => CLK, Q => 
                           REGISTERS_20_8_port, QN => n17265);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n3167, CK => CLK, Q => 
                           REGISTERS_20_7_port, QN => n17896);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n3166, CK => CLK, Q => 
                           REGISTERS_20_6_port, QN => n17897);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n3165, CK => CLK, Q => 
                           REGISTERS_20_5_port, QN => n17583);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n3164, CK => CLK, Q => 
                           REGISTERS_20_4_port, QN => n17584);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n3163, CK => CLK, Q => 
                           REGISTERS_20_3_port, QN => n17585);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n3162, CK => CLK, Q => 
                           REGISTERS_20_2_port, QN => n17898);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n3161, CK => CLK, Q => 
                           REGISTERS_20_1_port, QN => n17899);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n3160, CK => CLK, Q => 
                           REGISTERS_20_0_port, QN => n17900);
   REGISTERS_reg_21_63_inst : DFF_X1 port map( D => n3159, CK => CLK, Q => 
                           REGISTERS_21_63_port, QN => n18012);
   REGISTERS_reg_21_62_inst : DFF_X1 port map( D => n3158, CK => CLK, Q => 
                           REGISTERS_21_62_port, QN => n16895);
   REGISTERS_reg_21_61_inst : DFF_X1 port map( D => n3157, CK => CLK, Q => 
                           REGISTERS_21_61_port, QN => n16979);
   REGISTERS_reg_21_60_inst : DFF_X1 port map( D => n3156, CK => CLK, Q => 
                           REGISTERS_21_60_port, QN => n16896);
   REGISTERS_reg_21_59_inst : DFF_X1 port map( D => n3155, CK => CLK, Q => 
                           REGISTERS_21_59_port, QN => n16980);
   REGISTERS_reg_21_58_inst : DFF_X1 port map( D => n3154, CK => CLK, Q => 
                           REGISTERS_21_58_port, QN => n16981);
   REGISTERS_reg_21_57_inst : DFF_X1 port map( D => n3153, CK => CLK, Q => 
                           REGISTERS_21_57_port, QN => n16982);
   REGISTERS_reg_21_56_inst : DFF_X1 port map( D => n3152, CK => CLK, Q => 
                           REGISTERS_21_56_port, QN => n16983);
   REGISTERS_reg_21_55_inst : DFF_X1 port map( D => n3151, CK => CLK, Q => 
                           REGISTERS_21_55_port, QN => n16984);
   REGISTERS_reg_21_54_inst : DFF_X1 port map( D => n3150, CK => CLK, Q => 
                           REGISTERS_21_54_port, QN => n16897);
   REGISTERS_reg_21_53_inst : DFF_X1 port map( D => n3149, CK => CLK, Q => 
                           REGISTERS_21_53_port, QN => n16985);
   REGISTERS_reg_21_52_inst : DFF_X1 port map( D => n3148, CK => CLK, Q => 
                           REGISTERS_21_52_port, QN => n16898);
   REGISTERS_reg_21_51_inst : DFF_X1 port map( D => n3147, CK => CLK, Q => 
                           REGISTERS_21_51_port, QN => n17586);
   REGISTERS_reg_21_50_inst : DFF_X1 port map( D => n3146, CK => CLK, Q => 
                           REGISTERS_21_50_port, QN => n17266);
   REGISTERS_reg_21_49_inst : DFF_X1 port map( D => n3145, CK => CLK, Q => 
                           REGISTERS_21_49_port, QN => n17587);
   REGISTERS_reg_21_48_inst : DFF_X1 port map( D => n3144, CK => n13730, Q => 
                           REGISTERS_21_48_port, QN => n17267);
   REGISTERS_reg_21_47_inst : DFF_X1 port map( D => n3143, CK => CLK, Q => 
                           REGISTERS_21_47_port, QN => n17588);
   REGISTERS_reg_21_46_inst : DFF_X1 port map( D => n3142, CK => CLK, Q => 
                           REGISTERS_21_46_port, QN => n17589);
   REGISTERS_reg_21_45_inst : DFF_X1 port map( D => n3141, CK => CLK, Q => 
                           REGISTERS_21_45_port, QN => n17590);
   REGISTERS_reg_21_44_inst : DFF_X1 port map( D => n3140, CK => CLK, Q => 
                           REGISTERS_21_44_port, QN => n17591);
   REGISTERS_reg_21_43_inst : DFF_X1 port map( D => n3139, CK => CLK, Q => 
                           REGISTERS_21_43_port, QN => n17268);
   REGISTERS_reg_21_42_inst : DFF_X1 port map( D => n3138, CK => CLK, Q => 
                           REGISTERS_21_42_port, QN => n17592);
   REGISTERS_reg_21_41_inst : DFF_X1 port map( D => n3137, CK => CLK, Q => 
                           REGISTERS_21_41_port, QN => n17269);
   REGISTERS_reg_21_40_inst : DFF_X1 port map( D => n3136, CK => CLK, Q => 
                           REGISTERS_21_40_port, QN => n17593);
   REGISTERS_reg_21_39_inst : DFF_X1 port map( D => n3135, CK => CLK, Q => 
                           REGISTERS_21_39_port, QN => n17594);
   REGISTERS_reg_21_38_inst : DFF_X1 port map( D => n3134, CK => CLK, Q => 
                           REGISTERS_21_38_port, QN => n17270);
   REGISTERS_reg_21_37_inst : DFF_X1 port map( D => n3133, CK => CLK, Q => 
                           REGISTERS_21_37_port, QN => n17271);
   REGISTERS_reg_21_36_inst : DFF_X1 port map( D => n3132, CK => CLK, Q => 
                           REGISTERS_21_36_port, QN => n17272);
   REGISTERS_reg_21_35_inst : DFF_X1 port map( D => n3131, CK => CLK, Q => 
                           REGISTERS_21_35_port, QN => n17595);
   REGISTERS_reg_21_34_inst : DFF_X1 port map( D => n3130, CK => CLK, Q => 
                           REGISTERS_21_34_port, QN => n17596);
   REGISTERS_reg_21_33_inst : DFF_X1 port map( D => n3129, CK => CLK, Q => 
                           REGISTERS_21_33_port, QN => n17597);
   REGISTERS_reg_21_32_inst : DFF_X1 port map( D => n3128, CK => CLK, Q => 
                           REGISTERS_21_32_port, QN => n17598);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n3127, CK => CLK, Q => 
                           REGISTERS_21_31_port, QN => n17273);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n3126, CK => CLK, Q => 
                           REGISTERS_21_30_port, QN => n17274);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n3125, CK => CLK, Q => 
                           REGISTERS_21_29_port, QN => n17275);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n3124, CK => CLK, Q => 
                           REGISTERS_21_28_port, QN => n17276);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n3123, CK => CLK, Q => 
                           REGISTERS_21_27_port, QN => n16986);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n3122, CK => CLK, Q => 
                           REGISTERS_21_26_port, QN => n16899);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n3121, CK => CLK, Q => 
                           REGISTERS_21_25_port, QN => n16987);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n3120, CK => CLK, Q => 
                           REGISTERS_21_24_port, QN => n16900);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n3119, CK => CLK, Q => 
                           REGISTERS_21_23_port, QN => n16901);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n3118, CK => CLK, Q => 
                           REGISTERS_21_22_port, QN => n16902);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n3117, CK => CLK, Q => 
                           REGISTERS_21_21_port, QN => n16988);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n3116, CK => CLK, Q => 
                           REGISTERS_21_20_port, QN => n16903);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n3115, CK => CLK, Q => 
                           REGISTERS_21_19_port, QN => n16989);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n3114, CK => CLK, Q => 
                           REGISTERS_21_18_port, QN => n16990);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n3113, CK => CLK, Q => 
                           REGISTERS_21_17_port, QN => n16991);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n3112, CK => CLK, Q => 
                           REGISTERS_21_16_port, QN => n16904);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n3111, CK => CLK, Q => 
                           REGISTERS_21_15_port, QN => n17599);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n3110, CK => CLK, Q => 
                           REGISTERS_21_14_port, QN => n17600);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n3109, CK => CLK, Q => 
                           REGISTERS_21_13_port, QN => n17601);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n3108, CK => CLK, Q => 
                           REGISTERS_21_12_port, QN => n17602);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n3107, CK => CLK, Q => 
                           REGISTERS_21_11_port, QN => n17603);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n3106, CK => CLK, Q => 
                           REGISTERS_21_10_port, QN => n17604);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n3105, CK => CLK, Q => 
                           REGISTERS_21_9_port, QN => n17605);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n3104, CK => CLK, Q => 
                           REGISTERS_21_8_port, QN => n17277);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n3103, CK => CLK, Q => 
                           REGISTERS_21_7_port, QN => n17606);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n3102, CK => CLK, Q => 
                           REGISTERS_21_6_port, QN => n17607);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n3101, CK => CLK, Q => 
                           REGISTERS_21_5_port, QN => n17608);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n3100, CK => CLK, Q => 
                           REGISTERS_21_4_port, QN => n17278);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n3099, CK => CLK, Q => 
                           REGISTERS_21_3_port, QN => n17279);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n3098, CK => CLK, Q => 
                           REGISTERS_21_2_port, QN => n17609);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n3097, CK => CLK, Q => 
                           REGISTERS_21_1_port, QN => n17610);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n3096, CK => CLK, Q => 
                           REGISTERS_21_0_port, QN => n17611);
   REGISTERS_reg_22_63_inst : DFF_X1 port map( D => n3095, CK => CLK, Q => 
                           REGISTERS_22_63_port, QN => n18240);
   REGISTERS_reg_22_62_inst : DFF_X1 port map( D => n3094, CK => CLK, Q => 
                           REGISTERS_22_62_port, QN => n16905);
   REGISTERS_reg_22_61_inst : DFF_X1 port map( D => n3093, CK => CLK, Q => 
                           REGISTERS_22_61_port, QN => n16906);
   REGISTERS_reg_22_60_inst : DFF_X1 port map( D => n3092, CK => CLK, Q => 
                           REGISTERS_22_60_port, QN => n16992);
   REGISTERS_reg_22_59_inst : DFF_X1 port map( D => n3091, CK => CLK, Q => 
                           REGISTERS_22_59_port, QN => n16993);
   REGISTERS_reg_22_58_inst : DFF_X1 port map( D => n3090, CK => CLK, Q => 
                           REGISTERS_22_58_port, QN => n16994);
   REGISTERS_reg_22_57_inst : DFF_X1 port map( D => n3089, CK => CLK, Q => 
                           REGISTERS_22_57_port, QN => n16995);
   REGISTERS_reg_22_56_inst : DFF_X1 port map( D => n3088, CK => CLK, Q => 
                           REGISTERS_22_56_port, QN => n16996);
   REGISTERS_reg_22_55_inst : DFF_X1 port map( D => n3087, CK => CLK, Q => 
                           REGISTERS_22_55_port, QN => n16997);
   REGISTERS_reg_22_54_inst : DFF_X1 port map( D => n3086, CK => CLK, Q => 
                           REGISTERS_22_54_port, QN => n16907);
   REGISTERS_reg_22_53_inst : DFF_X1 port map( D => n3085, CK => CLK, Q => 
                           REGISTERS_22_53_port, QN => n17112);
   REGISTERS_reg_22_52_inst : DFF_X1 port map( D => n3084, CK => CLK, Q => 
                           REGISTERS_22_52_port, QN => n16998);
   REGISTERS_reg_22_51_inst : DFF_X1 port map( D => n3083, CK => CLK, Q => 
                           REGISTERS_22_51_port, QN => n17280);
   REGISTERS_reg_22_50_inst : DFF_X1 port map( D => n3082, CK => CLK, Q => 
                           REGISTERS_22_50_port, QN => n17281);
   REGISTERS_reg_22_49_inst : DFF_X1 port map( D => n3081, CK => CLK, Q => 
                           REGISTERS_22_49_port, QN => n17282);
   REGISTERS_reg_22_48_inst : DFF_X1 port map( D => n3080, CK => CLK, Q => 
                           REGISTERS_22_48_port, QN => n17283);
   REGISTERS_reg_22_47_inst : DFF_X1 port map( D => n3079, CK => CLK, Q => 
                           REGISTERS_22_47_port, QN => n17612);
   REGISTERS_reg_22_46_inst : DFF_X1 port map( D => n3078, CK => CLK, Q => 
                           REGISTERS_22_46_port, QN => n17284);
   REGISTERS_reg_22_45_inst : DFF_X1 port map( D => n3077, CK => CLK, Q => 
                           REGISTERS_22_45_port, QN => n17613);
   REGISTERS_reg_22_44_inst : DFF_X1 port map( D => n3076, CK => CLK, Q => 
                           REGISTERS_22_44_port, QN => n17285);
   REGISTERS_reg_22_43_inst : DFF_X1 port map( D => n3075, CK => CLK, Q => 
                           REGISTERS_22_43_port, QN => n17286);
   REGISTERS_reg_22_42_inst : DFF_X1 port map( D => n3074, CK => CLK, Q => 
                           REGISTERS_22_42_port, QN => n17614);
   REGISTERS_reg_22_41_inst : DFF_X1 port map( D => n3073, CK => CLK, Q => 
                           REGISTERS_22_41_port, QN => n17615);
   REGISTERS_reg_22_40_inst : DFF_X1 port map( D => n3072, CK => CLK, Q => 
                           REGISTERS_22_40_port, QN => n17616);
   REGISTERS_reg_22_39_inst : DFF_X1 port map( D => n3071, CK => CLK, Q => 
                           REGISTERS_22_39_port, QN => n17287);
   REGISTERS_reg_22_38_inst : DFF_X1 port map( D => n3070, CK => CLK, Q => 
                           REGISTERS_22_38_port, QN => n17288);
   REGISTERS_reg_22_37_inst : DFF_X1 port map( D => n3069, CK => CLK, Q => 
                           REGISTERS_22_37_port, QN => n17289);
   REGISTERS_reg_22_36_inst : DFF_X1 port map( D => n3068, CK => CLK, Q => 
                           REGISTERS_22_36_port, QN => n17617);
   REGISTERS_reg_22_35_inst : DFF_X1 port map( D => n3067, CK => CLK, Q => 
                           REGISTERS_22_35_port, QN => n17618);
   REGISTERS_reg_22_34_inst : DFF_X1 port map( D => n3066, CK => CLK, Q => 
                           REGISTERS_22_34_port, QN => n17290);
   REGISTERS_reg_22_33_inst : DFF_X1 port map( D => n3065, CK => CLK, Q => 
                           REGISTERS_22_33_port, QN => n17291);
   REGISTERS_reg_22_32_inst : DFF_X1 port map( D => n3064, CK => n13730, Q => 
                           REGISTERS_22_32_port, QN => n17619);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n3063, CK => CLK, Q => 
                           REGISTERS_22_31_port, QN => n17620);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n3062, CK => CLK, Q => 
                           REGISTERS_22_30_port, QN => n17621);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n3061, CK => CLK, Q => 
                           REGISTERS_22_29_port, QN => n17292);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n3060, CK => CLK, Q => 
                           REGISTERS_22_28_port, QN => n17622);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n3059, CK => CLK, Q => 
                           REGISTERS_22_27_port, QN => n16908);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n3058, CK => CLK, Q => 
                           REGISTERS_22_26_port, QN => n16909);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n3057, CK => CLK, Q => 
                           REGISTERS_22_25_port, QN => n16999);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n3056, CK => CLK, Q => 
                           REGISTERS_22_24_port, QN => n17000);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n3055, CK => CLK, Q => 
                           REGISTERS_22_23_port, QN => n16910);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n3054, CK => CLK, Q => 
                           REGISTERS_22_22_port, QN => n17001);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n3053, CK => CLK, Q => 
                           REGISTERS_22_21_port, QN => n16911);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n3052, CK => CLK, Q => 
                           REGISTERS_22_20_port, QN => n16912);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n3051, CK => CLK, Q => 
                           REGISTERS_22_19_port, QN => n17113);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n3050, CK => CLK, Q => 
                           REGISTERS_22_18_port, QN => n16913);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n3049, CK => CLK, Q => 
                           REGISTERS_22_17_port, QN => n16914);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n3048, CK => CLK, Q => 
                           REGISTERS_22_16_port, QN => n17002);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n3047, CK => CLK, Q => 
                           REGISTERS_22_15_port, QN => n17623);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n3046, CK => CLK, Q => 
                           REGISTERS_22_14_port, QN => n17293);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n3045, CK => CLK, Q => 
                           REGISTERS_22_13_port, QN => n17624);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n3044, CK => CLK, Q => 
                           REGISTERS_22_12_port, QN => n17294);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n3043, CK => CLK, Q => 
                           REGISTERS_22_11_port, QN => n17295);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n3042, CK => CLK, Q => 
                           REGISTERS_22_10_port, QN => n17625);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n3041, CK => CLK, Q => 
                           REGISTERS_22_9_port, QN => n17296);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n3040, CK => CLK, Q => 
                           REGISTERS_22_8_port, QN => n17297);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n3039, CK => CLK, Q => 
                           REGISTERS_22_7_port, QN => n17626);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n3038, CK => CLK, Q => 
                           REGISTERS_22_6_port, QN => n17298);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n3037, CK => CLK, Q => 
                           REGISTERS_22_5_port, QN => n17627);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n3036, CK => CLK, Q => 
                           REGISTERS_22_4_port, QN => n17299);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n3035, CK => CLK, Q => 
                           REGISTERS_22_3_port, QN => n17628);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n3034, CK => CLK, Q => 
                           REGISTERS_22_2_port, QN => n17300);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n3033, CK => CLK, Q => 
                           REGISTERS_22_1_port, QN => n17301);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n3032, CK => CLK, Q => 
                           REGISTERS_22_0_port, QN => n17629);
   REGISTERS_reg_23_63_inst : DFF_X1 port map( D => n3031, CK => CLK, Q => 
                           REGISTERS_23_63_port, QN => n18698);
   REGISTERS_reg_23_62_inst : DFF_X1 port map( D => n3030, CK => CLK, Q => 
                           REGISTERS_23_62_port, QN => n17003);
   REGISTERS_reg_23_61_inst : DFF_X1 port map( D => n3029, CK => CLK, Q => 
                           REGISTERS_23_61_port, QN => n17114);
   REGISTERS_reg_23_60_inst : DFF_X1 port map( D => n3028, CK => CLK, Q => 
                           REGISTERS_23_60_port, QN => n17004);
   REGISTERS_reg_23_59_inst : DFF_X1 port map( D => n3027, CK => CLK, Q => 
                           REGISTERS_23_59_port, QN => n17005);
   REGISTERS_reg_23_58_inst : DFF_X1 port map( D => n3026, CK => CLK, Q => 
                           REGISTERS_23_58_port, QN => n17006);
   REGISTERS_reg_23_57_inst : DFF_X1 port map( D => n3025, CK => CLK, Q => 
                           REGISTERS_23_57_port, QN => n17115);
   REGISTERS_reg_23_56_inst : DFF_X1 port map( D => n3024, CK => CLK, Q => 
                           REGISTERS_23_56_port, QN => n17007);
   REGISTERS_reg_23_55_inst : DFF_X1 port map( D => n3023, CK => CLK, Q => 
                           REGISTERS_23_55_port, QN => n16915);
   REGISTERS_reg_23_54_inst : DFF_X1 port map( D => n3022, CK => CLK, Q => 
                           REGISTERS_23_54_port, QN => n17008);
   REGISTERS_reg_23_53_inst : DFF_X1 port map( D => n3021, CK => CLK, Q => 
                           REGISTERS_23_53_port, QN => n17009);
   REGISTERS_reg_23_52_inst : DFF_X1 port map( D => n3020, CK => CLK, Q => 
                           REGISTERS_23_52_port, QN => n17116);
   REGISTERS_reg_23_51_inst : DFF_X1 port map( D => n3019, CK => CLK, Q => 
                           REGISTERS_23_51_port, QN => n17630);
   REGISTERS_reg_23_50_inst : DFF_X1 port map( D => n3018, CK => CLK, Q => 
                           REGISTERS_23_50_port, QN => n17631);
   REGISTERS_reg_23_49_inst : DFF_X1 port map( D => n3017, CK => CLK, Q => 
                           REGISTERS_23_49_port, QN => n17632);
   REGISTERS_reg_23_48_inst : DFF_X1 port map( D => n3016, CK => CLK, Q => 
                           REGISTERS_23_48_port, QN => n17633);
   REGISTERS_reg_23_47_inst : DFF_X1 port map( D => n3015, CK => CLK, Q => 
                           REGISTERS_23_47_port, QN => n17901);
   REGISTERS_reg_23_46_inst : DFF_X1 port map( D => n3014, CK => CLK, Q => 
                           REGISTERS_23_46_port, QN => n17902);
   REGISTERS_reg_23_45_inst : DFF_X1 port map( D => n3013, CK => CLK, Q => 
                           REGISTERS_23_45_port, QN => n17302);
   REGISTERS_reg_23_44_inst : DFF_X1 port map( D => n3012, CK => CLK, Q => 
                           REGISTERS_23_44_port, QN => n17634);
   REGISTERS_reg_23_43_inst : DFF_X1 port map( D => n3011, CK => CLK, Q => 
                           REGISTERS_23_43_port, QN => n17635);
   REGISTERS_reg_23_42_inst : DFF_X1 port map( D => n3010, CK => CLK, Q => 
                           REGISTERS_23_42_port, QN => n17903);
   REGISTERS_reg_23_41_inst : DFF_X1 port map( D => n3009, CK => CLK, Q => 
                           REGISTERS_23_41_port, QN => n17904);
   REGISTERS_reg_23_40_inst : DFF_X1 port map( D => n3008, CK => CLK, Q => 
                           REGISTERS_23_40_port, QN => n17303);
   REGISTERS_reg_23_39_inst : DFF_X1 port map( D => n3007, CK => CLK, Q => 
                           REGISTERS_23_39_port, QN => n17636);
   REGISTERS_reg_23_38_inst : DFF_X1 port map( D => n3006, CK => CLK, Q => 
                           REGISTERS_23_38_port, QN => n17637);
   REGISTERS_reg_23_37_inst : DFF_X1 port map( D => n3005, CK => CLK, Q => 
                           REGISTERS_23_37_port, QN => n17905);
   REGISTERS_reg_23_36_inst : DFF_X1 port map( D => n3004, CK => CLK, Q => 
                           REGISTERS_23_36_port, QN => n17906);
   REGISTERS_reg_23_35_inst : DFF_X1 port map( D => n3003, CK => CLK, Q => 
                           REGISTERS_23_35_port, QN => n17907);
   REGISTERS_reg_23_34_inst : DFF_X1 port map( D => n3002, CK => CLK, Q => 
                           REGISTERS_23_34_port, QN => n17304);
   REGISTERS_reg_23_33_inst : DFF_X1 port map( D => n3001, CK => CLK, Q => 
                           REGISTERS_23_33_port, QN => n17638);
   REGISTERS_reg_23_32_inst : DFF_X1 port map( D => n3000, CK => CLK, Q => 
                           REGISTERS_23_32_port, QN => n17305);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n2999, CK => CLK, Q => 
                           REGISTERS_23_31_port, QN => n17908);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n2998, CK => CLK, Q => 
                           REGISTERS_23_30_port, QN => n17909);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n2997, CK => CLK, Q => 
                           REGISTERS_23_29_port, QN => n17306);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n2996, CK => CLK, Q => 
                           REGISTERS_23_28_port, QN => n17639);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n2995, CK => CLK, Q => 
                           REGISTERS_23_27_port, QN => n17010);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n2994, CK => CLK, Q => 
                           REGISTERS_23_26_port, QN => n17011);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n2993, CK => CLK, Q => 
                           REGISTERS_23_25_port, QN => n16916);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n2992, CK => CLK, Q => 
                           REGISTERS_23_24_port, QN => n16917);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n2991, CK => CLK, Q => 
                           REGISTERS_23_23_port, QN => n16918);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n2990, CK => CLK, Q => 
                           REGISTERS_23_22_port, QN => n17117);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n2989, CK => CLK, Q => 
                           REGISTERS_23_21_port, QN => n17012);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n2988, CK => CLK, Q => 
                           REGISTERS_23_20_port, QN => n17118);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n2987, CK => CLK, Q => 
                           REGISTERS_23_19_port, QN => n17119);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n2986, CK => n13730, Q => 
                           REGISTERS_23_18_port, QN => n17013);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n2985, CK => CLK, Q => 
                           REGISTERS_23_17_port, QN => n17120);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n2984, CK => CLK, Q => 
                           REGISTERS_23_16_port, QN => n17014);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n2983, CK => CLK, Q => 
                           REGISTERS_23_15_port, QN => n17640);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n2982, CK => CLK, Q => 
                           REGISTERS_23_14_port, QN => n17641);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n2981, CK => CLK, Q => 
                           REGISTERS_23_13_port, QN => n17910);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n2980, CK => CLK, Q => 
                           REGISTERS_23_12_port, QN => n17642);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n2979, CK => CLK, Q => 
                           REGISTERS_23_11_port, QN => n17643);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n2978, CK => CLK, Q => 
                           REGISTERS_23_10_port, QN => n17644);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n2977, CK => CLK, Q => 
                           REGISTERS_23_9_port, QN => n17645);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n2976, CK => CLK, Q => 
                           REGISTERS_23_8_port, QN => n17307);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n2975, CK => CLK, Q => 
                           REGISTERS_23_7_port, QN => n17646);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n2974, CK => CLK, Q => 
                           REGISTERS_23_6_port, QN => n17911);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n2973, CK => CLK, Q => 
                           REGISTERS_23_5_port, QN => n17308);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n2972, CK => CLK, Q => 
                           REGISTERS_23_4_port, QN => n17647);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n2971, CK => CLK, Q => 
                           REGISTERS_23_3_port, QN => n17309);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n2970, CK => CLK, Q => 
                           REGISTERS_23_2_port, QN => n17310);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n2969, CK => CLK, Q => 
                           REGISTERS_23_1_port, QN => n17648);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n2968, CK => CLK, Q => 
                           REGISTERS_23_0_port, QN => n17649);
   REGISTERS_reg_24_63_inst : DFF_X1 port map( D => n2967, CK => CLK, Q => 
                           REGISTERS_24_63_port, QN => n18013);
   REGISTERS_reg_24_62_inst : DFF_X1 port map( D => n2966, CK => CLK, Q => 
                           REGISTERS_24_62_port, QN => n17015);
   REGISTERS_reg_24_61_inst : DFF_X1 port map( D => n2965, CK => CLK, Q => 
                           REGISTERS_24_61_port, QN => n17121);
   REGISTERS_reg_24_60_inst : DFF_X1 port map( D => n2964, CK => CLK, Q => 
                           REGISTERS_24_60_port, QN => n17122);
   REGISTERS_reg_24_59_inst : DFF_X1 port map( D => n2963, CK => CLK, Q => 
                           REGISTERS_24_59_port, QN => n17123);
   REGISTERS_reg_24_58_inst : DFF_X1 port map( D => n2962, CK => CLK, Q => 
                           REGISTERS_24_58_port, QN => n16919);
   REGISTERS_reg_24_57_inst : DFF_X1 port map( D => n2961, CK => CLK, Q => 
                           REGISTERS_24_57_port, QN => n17016);
   REGISTERS_reg_24_56_inst : DFF_X1 port map( D => n2960, CK => CLK, Q => 
                           REGISTERS_24_56_port, QN => n16920);
   REGISTERS_reg_24_55_inst : DFF_X1 port map( D => n2959, CK => CLK, Q => 
                           REGISTERS_24_55_port, QN => n17124);
   REGISTERS_reg_24_54_inst : DFF_X1 port map( D => n2958, CK => CLK, Q => 
                           REGISTERS_24_54_port, QN => n17125);
   REGISTERS_reg_24_53_inst : DFF_X1 port map( D => n2957, CK => CLK, Q => 
                           REGISTERS_24_53_port, QN => n16921);
   REGISTERS_reg_24_52_inst : DFF_X1 port map( D => n2956, CK => CLK, Q => 
                           REGISTERS_24_52_port, QN => n17017);
   REGISTERS_reg_24_51_inst : DFF_X1 port map( D => n2955, CK => CLK, Q => 
                           REGISTERS_24_51_port, QN => n17650);
   REGISTERS_reg_24_50_inst : DFF_X1 port map( D => n2954, CK => CLK, Q => 
                           REGISTERS_24_50_port, QN => n17651);
   REGISTERS_reg_24_49_inst : DFF_X1 port map( D => n2953, CK => CLK, Q => 
                           REGISTERS_24_49_port, QN => n17912);
   REGISTERS_reg_24_48_inst : DFF_X1 port map( D => n2952, CK => CLK, Q => 
                           REGISTERS_24_48_port, QN => n17652);
   REGISTERS_reg_24_47_inst : DFF_X1 port map( D => n2951, CK => CLK, Q => 
                           REGISTERS_24_47_port, QN => n17311);
   REGISTERS_reg_24_46_inst : DFF_X1 port map( D => n2950, CK => CLK, Q => 
                           REGISTERS_24_46_port, QN => n17653);
   REGISTERS_reg_24_45_inst : DFF_X1 port map( D => n2949, CK => CLK, Q => 
                           REGISTERS_24_45_port, QN => n17654);
   REGISTERS_reg_24_44_inst : DFF_X1 port map( D => n2948, CK => CLK, Q => 
                           REGISTERS_24_44_port, QN => n17312);
   REGISTERS_reg_24_43_inst : DFF_X1 port map( D => n2947, CK => CLK, Q => 
                           REGISTERS_24_43_port, QN => n17913);
   REGISTERS_reg_24_42_inst : DFF_X1 port map( D => n2946, CK => CLK, Q => 
                           REGISTERS_24_42_port, QN => n17313);
   REGISTERS_reg_24_41_inst : DFF_X1 port map( D => n2945, CK => CLK, Q => 
                           REGISTERS_24_41_port, QN => n17314);
   REGISTERS_reg_24_40_inst : DFF_X1 port map( D => n2944, CK => CLK, Q => 
                           REGISTERS_24_40_port, QN => n17655);
   REGISTERS_reg_24_39_inst : DFF_X1 port map( D => n2943, CK => CLK, Q => 
                           REGISTERS_24_39_port, QN => n17656);
   REGISTERS_reg_24_38_inst : DFF_X1 port map( D => n2942, CK => CLK, Q => 
                           REGISTERS_24_38_port, QN => n17914);
   REGISTERS_reg_24_37_inst : DFF_X1 port map( D => n2941, CK => CLK, Q => 
                           REGISTERS_24_37_port, QN => n17315);
   REGISTERS_reg_24_36_inst : DFF_X1 port map( D => n2940, CK => n13730, Q => 
                           REGISTERS_24_36_port, QN => n17316);
   REGISTERS_reg_24_35_inst : DFF_X1 port map( D => n2939, CK => CLK, Q => 
                           REGISTERS_24_35_port, QN => n17657);
   REGISTERS_reg_24_34_inst : DFF_X1 port map( D => n2938, CK => CLK, Q => 
                           REGISTERS_24_34_port, QN => n17915);
   REGISTERS_reg_24_33_inst : DFF_X1 port map( D => n2937, CK => CLK, Q => 
                           REGISTERS_24_33_port, QN => n17916);
   REGISTERS_reg_24_32_inst : DFF_X1 port map( D => n2936, CK => CLK, Q => 
                           REGISTERS_24_32_port, QN => n17917);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n2935, CK => CLK, Q => 
                           REGISTERS_24_31_port, QN => n17317);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n2934, CK => CLK, Q => 
                           REGISTERS_24_30_port, QN => n17318);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n2933, CK => CLK, Q => 
                           REGISTERS_24_29_port, QN => n17658);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n2932, CK => CLK, Q => 
                           REGISTERS_24_28_port, QN => n17319);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n2931, CK => CLK, Q => 
                           REGISTERS_24_27_port, QN => n17018);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n2930, CK => CLK, Q => 
                           REGISTERS_24_26_port, QN => n17019);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n2929, CK => CLK, Q => 
                           REGISTERS_24_25_port, QN => n17126);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n2928, CK => CLK, Q => 
                           REGISTERS_24_24_port, QN => n17127);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n2927, CK => CLK, Q => 
                           REGISTERS_24_23_port, QN => n17020);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n2926, CK => CLK, Q => 
                           REGISTERS_24_22_port, QN => n16922);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n2925, CK => CLK, Q => 
                           REGISTERS_24_21_port, QN => n17021);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n2924, CK => CLK, Q => 
                           REGISTERS_24_20_port, QN => n17022);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n2923, CK => CLK, Q => 
                           REGISTERS_24_19_port, QN => n16923);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n2922, CK => CLK, Q => 
                           REGISTERS_24_18_port, QN => n17023);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n2921, CK => CLK, Q => 
                           REGISTERS_24_17_port, QN => n17128);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n2920, CK => CLK, Q => 
                           REGISTERS_24_16_port, QN => n17024);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n2919, CK => CLK, Q => 
                           REGISTERS_24_15_port, QN => n17320);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n2918, CK => CLK, Q => 
                           REGISTERS_24_14_port, QN => n17918);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n2917, CK => CLK, Q => 
                           REGISTERS_24_13_port, QN => n17659);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n2916, CK => CLK, Q => 
                           REGISTERS_24_12_port, QN => n17660);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n2915, CK => CLK, Q => 
                           REGISTERS_24_11_port, QN => n17321);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n2914, CK => CLK, Q => 
                           REGISTERS_24_10_port, QN => n17919);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n2913, CK => CLK, Q => 
                           REGISTERS_24_9_port, QN => n17322);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n2912, CK => CLK, Q => 
                           REGISTERS_24_8_port, QN => n17920);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n2911, CK => CLK, Q => 
                           REGISTERS_24_7_port, QN => n17921);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n2910, CK => CLK, Q => 
                           REGISTERS_24_6_port, QN => n17661);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n2909, CK => CLK, Q => 
                           REGISTERS_24_5_port, QN => n17662);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n2908, CK => CLK, Q => 
                           REGISTERS_24_4_port, QN => n17323);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n2907, CK => CLK, Q => 
                           REGISTERS_24_3_port, QN => n17663);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n2906, CK => CLK, Q => 
                           REGISTERS_24_2_port, QN => n17922);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n2905, CK => CLK, Q => 
                           REGISTERS_24_1_port, QN => n17664);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n2904, CK => CLK, Q => 
                           REGISTERS_24_0_port, QN => n17665);
   REGISTERS_reg_25_63_inst : DFF_X1 port map( D => n2903, CK => CLK, Q => 
                           REGISTERS_25_63_port, QN => n18241);
   REGISTERS_reg_25_62_inst : DFF_X1 port map( D => n2902, CK => CLK, Q => 
                           REGISTERS_25_62_port, QN => n17025);
   REGISTERS_reg_25_61_inst : DFF_X1 port map( D => n2901, CK => CLK, Q => 
                           REGISTERS_25_61_port, QN => n16924);
   REGISTERS_reg_25_60_inst : DFF_X1 port map( D => n2900, CK => CLK, Q => 
                           REGISTERS_25_60_port, QN => n17129);
   REGISTERS_reg_25_59_inst : DFF_X1 port map( D => n2899, CK => CLK, Q => 
                           REGISTERS_25_59_port, QN => n17026);
   REGISTERS_reg_25_58_inst : DFF_X1 port map( D => n2898, CK => CLK, Q => 
                           REGISTERS_25_58_port, QN => n17130);
   REGISTERS_reg_25_57_inst : DFF_X1 port map( D => n2897, CK => CLK, Q => 
                           REGISTERS_25_57_port, QN => n17027);
   REGISTERS_reg_25_56_inst : DFF_X1 port map( D => n2896, CK => CLK, Q => 
                           REGISTERS_25_56_port, QN => n16925);
   REGISTERS_reg_25_55_inst : DFF_X1 port map( D => n2895, CK => CLK, Q => 
                           REGISTERS_25_55_port, QN => n17131);
   REGISTERS_reg_25_54_inst : DFF_X1 port map( D => n2894, CK => CLK, Q => 
                           REGISTERS_25_54_port, QN => n17132);
   REGISTERS_reg_25_53_inst : DFF_X1 port map( D => n2893, CK => CLK, Q => 
                           REGISTERS_25_53_port, QN => n17028);
   REGISTERS_reg_25_52_inst : DFF_X1 port map( D => n2892, CK => CLK, Q => 
                           REGISTERS_25_52_port, QN => n17029);
   REGISTERS_reg_25_51_inst : DFF_X1 port map( D => n2891, CK => CLK, Q => 
                           REGISTERS_25_51_port, QN => n17666);
   REGISTERS_reg_25_50_inst : DFF_X1 port map( D => n2890, CK => CLK, Q => 
                           REGISTERS_25_50_port, QN => n17923);
   REGISTERS_reg_25_49_inst : DFF_X1 port map( D => n2889, CK => CLK, Q => 
                           REGISTERS_25_49_port, QN => n17924);
   REGISTERS_reg_25_48_inst : DFF_X1 port map( D => n2888, CK => n13730, Q => 
                           REGISTERS_25_48_port, QN => n17925);
   REGISTERS_reg_25_47_inst : DFF_X1 port map( D => n2887, CK => CLK, Q => 
                           REGISTERS_25_47_port, QN => n17667);
   REGISTERS_reg_25_46_inst : DFF_X1 port map( D => n2886, CK => CLK, Q => 
                           REGISTERS_25_46_port, QN => n17926);
   REGISTERS_reg_25_45_inst : DFF_X1 port map( D => n2885, CK => CLK, Q => 
                           REGISTERS_25_45_port, QN => n17927);
   REGISTERS_reg_25_44_inst : DFF_X1 port map( D => n2884, CK => CLK, Q => 
                           REGISTERS_25_44_port, QN => n17928);
   REGISTERS_reg_25_43_inst : DFF_X1 port map( D => n2883, CK => n13730, Q => 
                           REGISTERS_25_43_port, QN => n17668);
   REGISTERS_reg_25_42_inst : DFF_X1 port map( D => n2882, CK => CLK, Q => 
                           REGISTERS_25_42_port, QN => n17669);
   REGISTERS_reg_25_41_inst : DFF_X1 port map( D => n2881, CK => CLK, Q => 
                           REGISTERS_25_41_port, QN => n17670);
   REGISTERS_reg_25_40_inst : DFF_X1 port map( D => n2880, CK => CLK, Q => 
                           REGISTERS_25_40_port, QN => n17671);
   REGISTERS_reg_25_39_inst : DFF_X1 port map( D => n2879, CK => CLK, Q => 
                           REGISTERS_25_39_port, QN => n17324);
   REGISTERS_reg_25_38_inst : DFF_X1 port map( D => n2878, CK => CLK, Q => 
                           REGISTERS_25_38_port, QN => n17929);
   REGISTERS_reg_25_37_inst : DFF_X1 port map( D => n2877, CK => CLK, Q => 
                           REGISTERS_25_37_port, QN => n17672);
   REGISTERS_reg_25_36_inst : DFF_X1 port map( D => n2876, CK => CLK, Q => 
                           REGISTERS_25_36_port, QN => n17930);
   REGISTERS_reg_25_35_inst : DFF_X1 port map( D => n2875, CK => CLK, Q => 
                           REGISTERS_25_35_port, QN => n17931);
   REGISTERS_reg_25_34_inst : DFF_X1 port map( D => n2874, CK => CLK, Q => 
                           REGISTERS_25_34_port, QN => n17673);
   REGISTERS_reg_25_33_inst : DFF_X1 port map( D => n2873, CK => CLK, Q => 
                           REGISTERS_25_33_port, QN => n17674);
   REGISTERS_reg_25_32_inst : DFF_X1 port map( D => n2872, CK => CLK, Q => 
                           REGISTERS_25_32_port, QN => n17675);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n2871, CK => CLK, Q => 
                           REGISTERS_25_31_port, QN => n17676);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n2870, CK => CLK, Q => 
                           REGISTERS_25_30_port, QN => n17932);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n2869, CK => CLK, Q => 
                           REGISTERS_25_29_port, QN => n17933);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n2868, CK => CLK, Q => 
                           REGISTERS_25_28_port, QN => n17934);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n2867, CK => CLK, Q => 
                           REGISTERS_25_27_port, QN => n17133);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n2866, CK => CLK, Q => 
                           REGISTERS_25_26_port, QN => n17134);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n2865, CK => CLK, Q => 
                           REGISTERS_25_25_port, QN => n17030);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n2864, CK => CLK, Q => 
                           REGISTERS_25_24_port, QN => n17031);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n2863, CK => CLK, Q => 
                           REGISTERS_25_23_port, QN => n17032);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n2862, CK => CLK, Q => 
                           REGISTERS_25_22_port, QN => n17033);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n2861, CK => CLK, Q => 
                           REGISTERS_25_21_port, QN => n17135);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n2860, CK => CLK, Q => 
                           REGISTERS_25_20_port, QN => n17136);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n2859, CK => CLK, Q => 
                           REGISTERS_25_19_port, QN => n16926);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n2858, CK => CLK, Q => 
                           REGISTERS_25_18_port, QN => n17034);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n2857, CK => CLK, Q => 
                           REGISTERS_25_17_port, QN => n17137);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n2856, CK => CLK, Q => 
                           REGISTERS_25_16_port, QN => n16927);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n2855, CK => CLK, Q => 
                           REGISTERS_25_15_port, QN => n17677);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n2854, CK => CLK, Q => 
                           REGISTERS_25_14_port, QN => n17678);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n2853, CK => CLK, Q => 
                           REGISTERS_25_13_port, QN => n17679);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n2852, CK => CLK, Q => 
                           REGISTERS_25_12_port, QN => n17680);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n2851, CK => CLK, Q => 
                           REGISTERS_25_11_port, QN => n17325);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n2850, CK => CLK, Q => 
                           REGISTERS_25_10_port, QN => n17681);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n2849, CK => CLK, Q => 
                           REGISTERS_25_9_port, QN => n17682);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n2848, CK => CLK, Q => 
                           REGISTERS_25_8_port, QN => n17683);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n2847, CK => CLK, Q => 
                           REGISTERS_25_7_port, QN => n17684);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n2846, CK => CLK, Q => 
                           REGISTERS_25_6_port, QN => n17935);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n2845, CK => CLK, Q => 
                           REGISTERS_25_5_port, QN => n17936);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n2844, CK => CLK, Q => 
                           REGISTERS_25_4_port, QN => n17937);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n2843, CK => CLK, Q => 
                           REGISTERS_25_3_port, QN => n17938);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n2842, CK => CLK, Q => 
                           REGISTERS_25_2_port, QN => n17939);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n2841, CK => CLK, Q => 
                           REGISTERS_25_1_port, QN => n17940);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n2840, CK => CLK, Q => 
                           REGISTERS_25_0_port, QN => n17685);
   REGISTERS_reg_26_63_inst : DFF_X1 port map( D => n2839, CK => CLK, Q => 
                           REGISTERS_26_63_port, QN => n18699);
   REGISTERS_reg_26_62_inst : DFF_X1 port map( D => n2838, CK => CLK, Q => 
                           REGISTERS_26_62_port, QN => n17138);
   REGISTERS_reg_26_61_inst : DFF_X1 port map( D => n2837, CK => CLK, Q => 
                           REGISTERS_26_61_port, QN => n17035);
   REGISTERS_reg_26_60_inst : DFF_X1 port map( D => n2836, CK => n13730, Q => 
                           REGISTERS_26_60_port, QN => n17036);
   REGISTERS_reg_26_59_inst : DFF_X1 port map( D => n2835, CK => CLK, Q => 
                           REGISTERS_26_59_port, QN => n17139);
   REGISTERS_reg_26_58_inst : DFF_X1 port map( D => n2834, CK => CLK, Q => 
                           REGISTERS_26_58_port, QN => n17037);
   REGISTERS_reg_26_57_inst : DFF_X1 port map( D => n2833, CK => CLK, Q => 
                           REGISTERS_26_57_port, QN => n17038);
   REGISTERS_reg_26_56_inst : DFF_X1 port map( D => n2832, CK => CLK, Q => 
                           REGISTERS_26_56_port, QN => n17140);
   REGISTERS_reg_26_55_inst : DFF_X1 port map( D => n2831, CK => n13730, Q => 
                           REGISTERS_26_55_port, QN => n17141);
   REGISTERS_reg_26_54_inst : DFF_X1 port map( D => n2830, CK => CLK, Q => 
                           REGISTERS_26_54_port, QN => n17039);
   REGISTERS_reg_26_53_inst : DFF_X1 port map( D => n2829, CK => CLK, Q => 
                           REGISTERS_26_53_port, QN => n17142);
   REGISTERS_reg_26_52_inst : DFF_X1 port map( D => n2828, CK => CLK, Q => 
                           REGISTERS_26_52_port, QN => n17143);
   REGISTERS_reg_26_51_inst : DFF_X1 port map( D => n2827, CK => CLK, Q => 
                           REGISTERS_26_51_port, QN => n17941);
   REGISTERS_reg_26_50_inst : DFF_X1 port map( D => n2826, CK => CLK, Q => 
                           REGISTERS_26_50_port, QN => n17942);
   REGISTERS_reg_26_49_inst : DFF_X1 port map( D => n2825, CK => CLK, Q => 
                           REGISTERS_26_49_port, QN => n17943);
   REGISTERS_reg_26_48_inst : DFF_X1 port map( D => n2824, CK => CLK, Q => 
                           REGISTERS_26_48_port, QN => n17686);
   REGISTERS_reg_26_47_inst : DFF_X1 port map( D => n2823, CK => CLK, Q => 
                           REGISTERS_26_47_port, QN => n17944);
   REGISTERS_reg_26_46_inst : DFF_X1 port map( D => n2822, CK => CLK, Q => 
                           REGISTERS_26_46_port, QN => n17687);
   REGISTERS_reg_26_45_inst : DFF_X1 port map( D => n2821, CK => CLK, Q => 
                           REGISTERS_26_45_port, QN => n17688);
   REGISTERS_reg_26_44_inst : DFF_X1 port map( D => n2820, CK => CLK, Q => 
                           REGISTERS_26_44_port, QN => n17945);
   REGISTERS_reg_26_43_inst : DFF_X1 port map( D => n2819, CK => CLK, Q => 
                           REGISTERS_26_43_port, QN => n17689);
   REGISTERS_reg_26_42_inst : DFF_X1 port map( D => n2818, CK => CLK, Q => 
                           REGISTERS_26_42_port, QN => n17946);
   REGISTERS_reg_26_41_inst : DFF_X1 port map( D => n2817, CK => CLK, Q => 
                           REGISTERS_26_41_port, QN => n17690);
   REGISTERS_reg_26_40_inst : DFF_X1 port map( D => n2816, CK => CLK, Q => 
                           REGISTERS_26_40_port, QN => n17691);
   REGISTERS_reg_26_39_inst : DFF_X1 port map( D => n2815, CK => CLK, Q => 
                           REGISTERS_26_39_port, QN => n17692);
   REGISTERS_reg_26_38_inst : DFF_X1 port map( D => n2814, CK => CLK, Q => 
                           REGISTERS_26_38_port, QN => n17947);
   REGISTERS_reg_26_37_inst : DFF_X1 port map( D => n2813, CK => CLK, Q => 
                           REGISTERS_26_37_port, QN => n17948);
   REGISTERS_reg_26_36_inst : DFF_X1 port map( D => n2812, CK => CLK, Q => 
                           REGISTERS_26_36_port, QN => n17949);
   REGISTERS_reg_26_35_inst : DFF_X1 port map( D => n2811, CK => CLK, Q => 
                           REGISTERS_26_35_port, QN => n17950);
   REGISTERS_reg_26_34_inst : DFF_X1 port map( D => n2810, CK => CLK, Q => 
                           REGISTERS_26_34_port, QN => n17951);
   REGISTERS_reg_26_33_inst : DFF_X1 port map( D => n2809, CK => CLK, Q => 
                           REGISTERS_26_33_port, QN => n17693);
   REGISTERS_reg_26_32_inst : DFF_X1 port map( D => n2808, CK => CLK, Q => 
                           REGISTERS_26_32_port, QN => n17694);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n2807, CK => CLK, Q => 
                           REGISTERS_26_31_port, QN => n17695);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n2806, CK => CLK, Q => 
                           REGISTERS_26_30_port, QN => n17696);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n2805, CK => CLK, Q => 
                           REGISTERS_26_29_port, QN => n17952);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n2804, CK => CLK, Q => 
                           REGISTERS_26_28_port, QN => n17953);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n2803, CK => CLK, Q => 
                           REGISTERS_26_27_port, QN => n17040);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n2802, CK => CLK, Q => 
                           REGISTERS_26_26_port, QN => n17144);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n2801, CK => CLK, Q => 
                           REGISTERS_26_25_port, QN => n17145);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n2800, CK => CLK, Q => 
                           REGISTERS_26_24_port, QN => n17041);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n2799, CK => CLK, Q => 
                           REGISTERS_26_23_port, QN => n17042);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n2798, CK => CLK, Q => 
                           REGISTERS_26_22_port, QN => n17146);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n2797, CK => CLK, Q => 
                           REGISTERS_26_21_port, QN => n17147);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n2796, CK => CLK, Q => 
                           REGISTERS_26_20_port, QN => n17043);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n2795, CK => CLK, Q => 
                           REGISTERS_26_19_port, QN => n17044);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n2794, CK => CLK, Q => 
                           REGISTERS_26_18_port, QN => n17045);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n2793, CK => CLK, Q => 
                           REGISTERS_26_17_port, QN => n17148);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n2792, CK => CLK, Q => 
                           REGISTERS_26_16_port, QN => n17149);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n2791, CK => CLK, Q => 
                           REGISTERS_26_15_port, QN => n17954);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n2790, CK => CLK, Q => 
                           REGISTERS_26_14_port, QN => n17955);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n2789, CK => CLK, Q => 
                           REGISTERS_26_13_port, QN => n17956);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n2788, CK => CLK, Q => 
                           REGISTERS_26_12_port, QN => n17697);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n2787, CK => CLK, Q => 
                           REGISTERS_26_11_port, QN => n17957);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n2786, CK => CLK, Q => 
                           REGISTERS_26_10_port, QN => n17698);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n2785, CK => CLK, Q => 
                           REGISTERS_26_9_port, QN => n17958);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n2784, CK => CLK, Q => 
                           REGISTERS_26_8_port, QN => n17959);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n2783, CK => CLK, Q => 
                           REGISTERS_26_7_port, QN => n17699);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n2782, CK => CLK, Q => 
                           REGISTERS_26_6_port, QN => n17700);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n2781, CK => CLK, Q => 
                           REGISTERS_26_5_port, QN => n17701);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n2780, CK => CLK, Q => 
                           REGISTERS_26_4_port, QN => n17960);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n2779, CK => CLK, Q => 
                           REGISTERS_26_3_port, QN => n17961);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n2778, CK => CLK, Q => 
                           REGISTERS_26_2_port, QN => n17962);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n2777, CK => CLK, Q => 
                           REGISTERS_26_1_port, QN => n17702);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n2776, CK => CLK, Q => 
                           REGISTERS_26_0_port, QN => n17703);
   REGISTERS_reg_27_63_inst : DFF_X1 port map( D => n2775, CK => CLK, Q => 
                           REGISTERS_27_63_port, QN => n18014);
   REGISTERS_reg_27_62_inst : DFF_X1 port map( D => n2774, CK => CLK, Q => 
                           REGISTERS_27_62_port, QN => n17150);
   REGISTERS_reg_27_61_inst : DFF_X1 port map( D => n2773, CK => CLK, Q => 
                           REGISTERS_27_61_port, QN => n16928);
   REGISTERS_reg_27_60_inst : DFF_X1 port map( D => n2772, CK => CLK, Q => 
                           REGISTERS_27_60_port, QN => n17046);
   REGISTERS_reg_27_59_inst : DFF_X1 port map( D => n2771, CK => CLK, Q => 
                           REGISTERS_27_59_port, QN => n17151);
   REGISTERS_reg_27_58_inst : DFF_X1 port map( D => n2770, CK => CLK, Q => 
                           REGISTERS_27_58_port, QN => n17047);
   REGISTERS_reg_27_57_inst : DFF_X1 port map( D => n2769, CK => CLK, Q => 
                           REGISTERS_27_57_port, QN => n16929);
   REGISTERS_reg_27_56_inst : DFF_X1 port map( D => n2768, CK => n13730, Q => 
                           REGISTERS_27_56_port, QN => n17152);
   REGISTERS_reg_27_55_inst : DFF_X1 port map( D => n2767, CK => CLK, Q => 
                           REGISTERS_27_55_port, QN => n16930);
   REGISTERS_reg_27_54_inst : DFF_X1 port map( D => n2766, CK => CLK, Q => 
                           REGISTERS_27_54_port, QN => n17048);
   REGISTERS_reg_27_53_inst : DFF_X1 port map( D => n2765, CK => CLK, Q => 
                           REGISTERS_27_53_port, QN => n17049);
   REGISTERS_reg_27_52_inst : DFF_X1 port map( D => n2764, CK => CLK, Q => 
                           REGISTERS_27_52_port, QN => n17050);
   REGISTERS_reg_27_51_inst : DFF_X1 port map( D => n2763, CK => CLK, Q => 
                           REGISTERS_27_51_port, QN => n17326);
   REGISTERS_reg_27_50_inst : DFF_X1 port map( D => n2762, CK => CLK, Q => 
                           REGISTERS_27_50_port, QN => n17963);
   REGISTERS_reg_27_49_inst : DFF_X1 port map( D => n2761, CK => CLK, Q => 
                           REGISTERS_27_49_port, QN => n17704);
   REGISTERS_reg_27_48_inst : DFF_X1 port map( D => n2760, CK => CLK, Q => 
                           REGISTERS_27_48_port, QN => n17705);
   REGISTERS_reg_27_47_inst : DFF_X1 port map( D => n2759, CK => CLK, Q => 
                           REGISTERS_27_47_port, QN => n17964);
   REGISTERS_reg_27_46_inst : DFF_X1 port map( D => n2758, CK => CLK, Q => 
                           REGISTERS_27_46_port, QN => n17706);
   REGISTERS_reg_27_45_inst : DFF_X1 port map( D => n2757, CK => CLK, Q => 
                           REGISTERS_27_45_port, QN => n17327);
   REGISTERS_reg_27_44_inst : DFF_X1 port map( D => n2756, CK => CLK, Q => 
                           REGISTERS_27_44_port, QN => n17965);
   REGISTERS_reg_27_43_inst : DFF_X1 port map( D => n2755, CK => CLK, Q => 
                           REGISTERS_27_43_port, QN => n17328);
   REGISTERS_reg_27_42_inst : DFF_X1 port map( D => n2754, CK => CLK, Q => 
                           REGISTERS_27_42_port, QN => n17707);
   REGISTERS_reg_27_41_inst : DFF_X1 port map( D => n2753, CK => CLK, Q => 
                           REGISTERS_27_41_port, QN => n17966);
   REGISTERS_reg_27_40_inst : DFF_X1 port map( D => n2752, CK => CLK, Q => 
                           REGISTERS_27_40_port, QN => n17967);
   REGISTERS_reg_27_39_inst : DFF_X1 port map( D => n2751, CK => CLK, Q => 
                           REGISTERS_27_39_port, QN => n17968);
   REGISTERS_reg_27_38_inst : DFF_X1 port map( D => n2750, CK => CLK, Q => 
                           REGISTERS_27_38_port, QN => n17708);
   REGISTERS_reg_27_37_inst : DFF_X1 port map( D => n2749, CK => CLK, Q => 
                           REGISTERS_27_37_port, QN => n17969);
   REGISTERS_reg_27_36_inst : DFF_X1 port map( D => n2748, CK => CLK, Q => 
                           REGISTERS_27_36_port, QN => n17709);
   REGISTERS_reg_27_35_inst : DFF_X1 port map( D => n2747, CK => n13730, Q => 
                           REGISTERS_27_35_port, QN => n17970);
   REGISTERS_reg_27_34_inst : DFF_X1 port map( D => n2746, CK => CLK, Q => 
                           REGISTERS_27_34_port, QN => n17710);
   REGISTERS_reg_27_33_inst : DFF_X1 port map( D => n2745, CK => CLK, Q => 
                           REGISTERS_27_33_port, QN => n17711);
   REGISTERS_reg_27_32_inst : DFF_X1 port map( D => n2744, CK => CLK, Q => 
                           REGISTERS_27_32_port, QN => n17971);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n2743, CK => CLK, Q => 
                           REGISTERS_27_31_port, QN => n17972);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n2742, CK => CLK, Q => 
                           REGISTERS_27_30_port, QN => n17712);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n2741, CK => CLK, Q => 
                           REGISTERS_27_29_port, QN => n17713);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n2740, CK => CLK, Q => 
                           REGISTERS_27_28_port, QN => n17714);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n2739, CK => CLK, Q => 
                           REGISTERS_27_27_port, QN => n17153);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n2738, CK => CLK, Q => 
                           REGISTERS_27_26_port, QN => n17154);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n2737, CK => CLK, Q => 
                           REGISTERS_27_25_port, QN => n17155);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n2736, CK => CLK, Q => 
                           REGISTERS_27_24_port, QN => n17156);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n2735, CK => CLK, Q => 
                           REGISTERS_27_23_port, QN => n17051);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n2734, CK => CLK, Q => 
                           REGISTERS_27_22_port, QN => n17052);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n2733, CK => CLK, Q => 
                           REGISTERS_27_21_port, QN => n16931);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n2732, CK => CLK, Q => 
                           REGISTERS_27_20_port, QN => n17053);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n2731, CK => CLK, Q => 
                           REGISTERS_27_19_port, QN => n17157);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n2730, CK => CLK, Q => 
                           REGISTERS_27_18_port, QN => n17158);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n2729, CK => CLK, Q => 
                           REGISTERS_27_17_port, QN => n17054);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n2728, CK => CLK, Q => 
                           REGISTERS_27_16_port, QN => n16932);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n2727, CK => CLK, Q => 
                           REGISTERS_27_15_port, QN => n17973);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n2726, CK => CLK, Q => 
                           REGISTERS_27_14_port, QN => n17329);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n2725, CK => n13730, Q => 
                           REGISTERS_27_13_port, QN => n17715);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n2724, CK => CLK, Q => 
                           REGISTERS_27_12_port, QN => n17974);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n2723, CK => CLK, Q => 
                           REGISTERS_27_11_port, QN => n17716);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n2722, CK => CLK, Q => 
                           REGISTERS_27_10_port, QN => n17975);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n2721, CK => CLK, Q => 
                           REGISTERS_27_9_port, QN => n17717);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n2720, CK => CLK, Q => 
                           REGISTERS_27_8_port, QN => n17718);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n2719, CK => CLK, Q => 
                           REGISTERS_27_7_port, QN => n17976);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n2718, CK => CLK, Q => 
                           REGISTERS_27_6_port, QN => n17977);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n2717, CK => CLK, Q => 
                           REGISTERS_27_5_port, QN => n17719);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n2716, CK => CLK, Q => 
                           REGISTERS_27_4_port, QN => n17720);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n2715, CK => CLK, Q => 
                           REGISTERS_27_3_port, QN => n17721);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n2714, CK => CLK, Q => 
                           REGISTERS_27_2_port, QN => n17330);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n2713, CK => CLK, Q => 
                           REGISTERS_27_1_port, QN => n17978);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n2712, CK => CLK, Q => 
                           REGISTERS_27_0_port, QN => n17722);
   REGISTERS_reg_28_63_inst : DFF_X1 port map( D => n2711, CK => CLK, Q => 
                           REGISTERS_28_63_port, QN => n18700);
   REGISTERS_reg_28_62_inst : DFF_X1 port map( D => n2710, CK => CLK, Q => 
                           REGISTERS_28_62_port, QN => n16933);
   REGISTERS_reg_28_61_inst : DFF_X1 port map( D => n2709, CK => CLK, Q => 
                           REGISTERS_28_61_port, QN => n17055);
   REGISTERS_reg_28_60_inst : DFF_X1 port map( D => n2708, CK => CLK, Q => 
                           REGISTERS_28_60_port, QN => n16934);
   REGISTERS_reg_28_59_inst : DFF_X1 port map( D => n2707, CK => CLK, Q => 
                           REGISTERS_28_59_port, QN => n17056);
   REGISTERS_reg_28_58_inst : DFF_X1 port map( D => n2706, CK => CLK, Q => 
                           REGISTERS_28_58_port, QN => n17057);
   REGISTERS_reg_28_57_inst : DFF_X1 port map( D => n2705, CK => CLK, Q => 
                           REGISTERS_28_57_port, QN => n17058);
   REGISTERS_reg_28_56_inst : DFF_X1 port map( D => n2704, CK => CLK, Q => 
                           REGISTERS_28_56_port, QN => n17059);
   REGISTERS_reg_28_55_inst : DFF_X1 port map( D => n2703, CK => CLK, Q => 
                           REGISTERS_28_55_port, QN => n17060);
   REGISTERS_reg_28_54_inst : DFF_X1 port map( D => n2702, CK => CLK, Q => 
                           REGISTERS_28_54_port, QN => n17061);
   REGISTERS_reg_28_53_inst : DFF_X1 port map( D => n2701, CK => CLK, Q => 
                           REGISTERS_28_53_port, QN => n17062);
   REGISTERS_reg_28_52_inst : DFF_X1 port map( D => n2700, CK => CLK, Q => 
                           REGISTERS_28_52_port, QN => n16935);
   REGISTERS_reg_28_51_inst : DFF_X1 port map( D => n2699, CK => CLK, Q => 
                           REGISTERS_28_51_port, QN => n17723);
   REGISTERS_reg_28_50_inst : DFF_X1 port map( D => n2698, CK => CLK, Q => 
                           REGISTERS_28_50_port, QN => n17724);
   REGISTERS_reg_28_49_inst : DFF_X1 port map( D => n2697, CK => CLK, Q => 
                           REGISTERS_28_49_port, QN => n17725);
   REGISTERS_reg_28_48_inst : DFF_X1 port map( D => n2696, CK => CLK, Q => 
                           REGISTERS_28_48_port, QN => n17979);
   REGISTERS_reg_28_47_inst : DFF_X1 port map( D => n2695, CK => CLK, Q => 
                           REGISTERS_28_47_port, QN => n17331);
   REGISTERS_reg_28_46_inst : DFF_X1 port map( D => n2694, CK => CLK, Q => 
                           REGISTERS_28_46_port, QN => n17726);
   REGISTERS_reg_28_45_inst : DFF_X1 port map( D => n2693, CK => CLK, Q => 
                           REGISTERS_28_45_port, QN => n17727);
   REGISTERS_reg_28_44_inst : DFF_X1 port map( D => n2692, CK => CLK, Q => 
                           REGISTERS_28_44_port, QN => n17728);
   REGISTERS_reg_28_43_inst : DFF_X1 port map( D => n2691, CK => CLK, Q => 
                           REGISTERS_28_43_port, QN => n17729);
   REGISTERS_reg_28_42_inst : DFF_X1 port map( D => n2690, CK => CLK, Q => 
                           REGISTERS_28_42_port, QN => n17332);
   REGISTERS_reg_28_41_inst : DFF_X1 port map( D => n2689, CK => CLK, Q => 
                           REGISTERS_28_41_port, QN => n17333);
   REGISTERS_reg_28_40_inst : DFF_X1 port map( D => n2688, CK => CLK, Q => 
                           REGISTERS_28_40_port, QN => n17334);
   REGISTERS_reg_28_39_inst : DFF_X1 port map( D => n2687, CK => CLK, Q => 
                           REGISTERS_28_39_port, QN => n17335);
   REGISTERS_reg_28_38_inst : DFF_X1 port map( D => n2686, CK => CLK, Q => 
                           REGISTERS_28_38_port, QN => n17730);
   REGISTERS_reg_28_37_inst : DFF_X1 port map( D => n2685, CK => CLK, Q => 
                           REGISTERS_28_37_port, QN => n17731);
   REGISTERS_reg_28_36_inst : DFF_X1 port map( D => n2684, CK => n13730, Q => 
                           REGISTERS_28_36_port, QN => n17732);
   REGISTERS_reg_28_35_inst : DFF_X1 port map( D => n2683, CK => CLK, Q => 
                           REGISTERS_28_35_port, QN => n17336);
   REGISTERS_reg_28_34_inst : DFF_X1 port map( D => n2682, CK => CLK, Q => 
                           REGISTERS_28_34_port, QN => n17733);
   REGISTERS_reg_28_33_inst : DFF_X1 port map( D => n2681, CK => CLK, Q => 
                           REGISTERS_28_33_port, QN => n17734);
   REGISTERS_reg_28_32_inst : DFF_X1 port map( D => n2680, CK => CLK, Q => 
                           REGISTERS_28_32_port, QN => n17735);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n2679, CK => CLK, Q => 
                           REGISTERS_28_31_port, QN => n17736);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n2678, CK => CLK, Q => 
                           REGISTERS_28_30_port, QN => n17980);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n2677, CK => CLK, Q => 
                           REGISTERS_28_29_port, QN => n17337);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n2676, CK => CLK, Q => 
                           REGISTERS_28_28_port, QN => n17737);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n2675, CK => CLK, Q => 
                           REGISTERS_28_27_port, QN => n17063);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n2674, CK => CLK, Q => 
                           REGISTERS_28_26_port, QN => n16936);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n2673, CK => CLK, Q => 
                           REGISTERS_28_25_port, QN => n16937);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n2672, CK => CLK, Q => 
                           REGISTERS_28_24_port, QN => n17064);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n2671, CK => CLK, Q => 
                           REGISTERS_28_23_port, QN => n16938);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n2670, CK => CLK, Q => 
                           REGISTERS_28_22_port, QN => n17065);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n2669, CK => CLK, Q => 
                           REGISTERS_28_21_port, QN => n16939);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n2668, CK => CLK, Q => 
                           REGISTERS_28_20_port, QN => n17066);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n2667, CK => CLK, Q => 
                           REGISTERS_28_19_port, QN => n17067);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n2666, CK => CLK, Q => 
                           REGISTERS_28_18_port, QN => n16940);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n2665, CK => CLK, Q => 
                           REGISTERS_28_17_port, QN => n16941);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n2664, CK => CLK, Q => 
                           REGISTERS_28_16_port, QN => n17068);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n2663, CK => CLK, Q => 
                           REGISTERS_28_15_port, QN => n17981);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n2662, CK => CLK, Q => 
                           REGISTERS_28_14_port, QN => n17338);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n2661, CK => CLK, Q => 
                           REGISTERS_28_13_port, QN => n17738);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n2660, CK => CLK, Q => 
                           REGISTERS_28_12_port, QN => n17739);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n2659, CK => CLK, Q => 
                           REGISTERS_28_11_port, QN => n17339);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n2658, CK => CLK, Q => 
                           REGISTERS_28_10_port, QN => n17340);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n2657, CK => CLK, Q => 
                           REGISTERS_28_9_port, QN => n17740);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n2656, CK => CLK, Q => 
                           REGISTERS_28_8_port, QN => n17741);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n2655, CK => CLK, Q => 
                           REGISTERS_28_7_port, QN => n17341);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n2654, CK => CLK, Q => 
                           REGISTERS_28_6_port, QN => n17742);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n2653, CK => CLK, Q => 
                           REGISTERS_28_5_port, QN => n17743);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n2652, CK => CLK, Q => 
                           REGISTERS_28_4_port, QN => n17744);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n2651, CK => CLK, Q => 
                           REGISTERS_28_3_port, QN => n17745);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n2650, CK => CLK, Q => 
                           REGISTERS_28_2_port, QN => n17746);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n2649, CK => CLK, Q => 
                           REGISTERS_28_1_port, QN => n17342);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n2648, CK => CLK, Q => 
                           REGISTERS_28_0_port, QN => n17982);
   REGISTERS_reg_29_63_inst : DFF_X1 port map( D => n2647, CK => CLK, Q => 
                           REGISTERS_29_63_port, QN => n18015);
   REGISTERS_reg_29_62_inst : DFF_X1 port map( D => n2646, CK => CLK, Q => 
                           REGISTERS_29_62_port, QN => n17069);
   REGISTERS_reg_29_61_inst : DFF_X1 port map( D => n2645, CK => CLK, Q => 
                           REGISTERS_29_61_port, QN => n17070);
   REGISTERS_reg_29_60_inst : DFF_X1 port map( D => n2644, CK => CLK, Q => 
                           REGISTERS_29_60_port, QN => n17071);
   REGISTERS_reg_29_59_inst : DFF_X1 port map( D => n2643, CK => CLK, Q => 
                           REGISTERS_29_59_port, QN => n16942);
   REGISTERS_reg_29_58_inst : DFF_X1 port map( D => n2642, CK => CLK, Q => 
                           REGISTERS_29_58_port, QN => n17072);
   REGISTERS_reg_29_57_inst : DFF_X1 port map( D => n2641, CK => CLK, Q => 
                           REGISTERS_29_57_port, QN => n16943);
   REGISTERS_reg_29_56_inst : DFF_X1 port map( D => n2640, CK => CLK, Q => 
                           REGISTERS_29_56_port, QN => n16944);
   REGISTERS_reg_29_55_inst : DFF_X1 port map( D => n2639, CK => CLK, Q => 
                           REGISTERS_29_55_port, QN => n16945);
   REGISTERS_reg_29_54_inst : DFF_X1 port map( D => n2638, CK => CLK, Q => 
                           REGISTERS_29_54_port, QN => n16946);
   REGISTERS_reg_29_53_inst : DFF_X1 port map( D => n2637, CK => CLK, Q => 
                           REGISTERS_29_53_port, QN => n16947);
   REGISTERS_reg_29_52_inst : DFF_X1 port map( D => n2636, CK => CLK, Q => 
                           REGISTERS_29_52_port, QN => n16948);
   REGISTERS_reg_29_51_inst : DFF_X1 port map( D => n2635, CK => CLK, Q => 
                           REGISTERS_29_51_port, QN => n17747);
   REGISTERS_reg_29_50_inst : DFF_X1 port map( D => n2634, CK => CLK, Q => 
                           REGISTERS_29_50_port, QN => n17343);
   REGISTERS_reg_29_49_inst : DFF_X1 port map( D => n2633, CK => CLK, Q => 
                           REGISTERS_29_49_port, QN => n17344);
   REGISTERS_reg_29_48_inst : DFF_X1 port map( D => n2632, CK => CLK, Q => 
                           REGISTERS_29_48_port, QN => n17345);
   REGISTERS_reg_29_47_inst : DFF_X1 port map( D => n2631, CK => CLK, Q => 
                           REGISTERS_29_47_port, QN => n17346);
   REGISTERS_reg_29_46_inst : DFF_X1 port map( D => n2630, CK => CLK, Q => 
                           REGISTERS_29_46_port, QN => n17347);
   REGISTERS_reg_29_45_inst : DFF_X1 port map( D => n2629, CK => CLK, Q => 
                           REGISTERS_29_45_port, QN => n17748);
   REGISTERS_reg_29_44_inst : DFF_X1 port map( D => n2628, CK => CLK, Q => 
                           REGISTERS_29_44_port, QN => n17348);
   REGISTERS_reg_29_43_inst : DFF_X1 port map( D => n2627, CK => CLK, Q => 
                           REGISTERS_29_43_port, QN => n17349);
   REGISTERS_reg_29_42_inst : DFF_X1 port map( D => n2626, CK => CLK, Q => 
                           REGISTERS_29_42_port, QN => n17350);
   REGISTERS_reg_29_41_inst : DFF_X1 port map( D => n2625, CK => CLK, Q => 
                           REGISTERS_29_41_port, QN => n17351);
   REGISTERS_reg_29_40_inst : DFF_X1 port map( D => n2624, CK => CLK, Q => 
                           REGISTERS_29_40_port, QN => n17983);
   REGISTERS_reg_29_39_inst : DFF_X1 port map( D => n2623, CK => CLK, Q => 
                           REGISTERS_29_39_port, QN => n17749);
   REGISTERS_reg_29_38_inst : DFF_X1 port map( D => n2622, CK => CLK, Q => 
                           REGISTERS_29_38_port, QN => n17750);
   REGISTERS_reg_29_37_inst : DFF_X1 port map( D => n2621, CK => CLK, Q => 
                           REGISTERS_29_37_port, QN => n17751);
   REGISTERS_reg_29_36_inst : DFF_X1 port map( D => n2620, CK => CLK, Q => 
                           REGISTERS_29_36_port, QN => n17984);
   REGISTERS_reg_29_35_inst : DFF_X1 port map( D => n2619, CK => CLK, Q => 
                           REGISTERS_29_35_port, QN => n17985);
   REGISTERS_reg_29_34_inst : DFF_X1 port map( D => n2618, CK => CLK, Q => 
                           REGISTERS_29_34_port, QN => n17752);
   REGISTERS_reg_29_33_inst : DFF_X1 port map( D => n2617, CK => CLK, Q => 
                           REGISTERS_29_33_port, QN => n17753);
   REGISTERS_reg_29_32_inst : DFF_X1 port map( D => n2616, CK => CLK, Q => 
                           REGISTERS_29_32_port, QN => n17352);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n2615, CK => CLK, Q => 
                           REGISTERS_29_31_port, QN => n17754);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n2614, CK => CLK, Q => 
                           REGISTERS_29_30_port, QN => n17353);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n2613, CK => CLK, Q => 
                           REGISTERS_29_29_port, QN => n17755);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n2612, CK => CLK, Q => 
                           REGISTERS_29_28_port, QN => n17354);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n2611, CK => CLK, Q => 
                           REGISTERS_29_27_port, QN => n17073);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n2610, CK => CLK, Q => 
                           REGISTERS_29_26_port, QN => n17074);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n2609, CK => CLK, Q => 
                           REGISTERS_29_25_port, QN => n16949);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n2608, CK => CLK, Q => 
                           REGISTERS_29_24_port, QN => n17075);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n2607, CK => n13730, Q => 
                           REGISTERS_29_23_port, QN => n16950);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n2606, CK => CLK, Q => 
                           REGISTERS_29_22_port, QN => n17076);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n2605, CK => CLK, Q => 
                           REGISTERS_29_21_port, QN => n17077);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n2604, CK => CLK, Q => 
                           REGISTERS_29_20_port, QN => n17078);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n2603, CK => CLK, Q => 
                           REGISTERS_29_19_port, QN => n16951);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n2602, CK => CLK, Q => 
                           REGISTERS_29_18_port, QN => n17079);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n2601, CK => CLK, Q => 
                           REGISTERS_29_17_port, QN => n16952);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n2600, CK => CLK, Q => 
                           REGISTERS_29_16_port, QN => n16953);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n2599, CK => CLK, Q => 
                           REGISTERS_29_15_port, QN => n17986);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n2598, CK => CLK, Q => 
                           REGISTERS_29_14_port, QN => n17756);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n2597, CK => CLK, Q => 
                           REGISTERS_29_13_port, QN => n17355);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n2596, CK => CLK, Q => 
                           REGISTERS_29_12_port, QN => n17356);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n2595, CK => CLK, Q => 
                           REGISTERS_29_11_port, QN => n17357);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n2594, CK => CLK, Q => 
                           REGISTERS_29_10_port, QN => n17987);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n2593, CK => CLK, Q => 
                           REGISTERS_29_9_port, QN => n17757);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n2592, CK => CLK, Q => 
                           REGISTERS_29_8_port, QN => n17988);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n2591, CK => CLK, Q => 
                           REGISTERS_29_7_port, QN => n17358);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n2590, CK => CLK, Q => 
                           REGISTERS_29_6_port, QN => n17359);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n2589, CK => CLK, Q => 
                           REGISTERS_29_5_port, QN => n17360);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n2588, CK => CLK, Q => 
                           REGISTERS_29_4_port, QN => n17361);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n2587, CK => CLK, Q => 
                           REGISTERS_29_3_port, QN => n17362);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n2586, CK => CLK, Q => 
                           REGISTERS_29_2_port, QN => n17363);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n2585, CK => CLK, Q => 
                           REGISTERS_29_1_port, QN => n17758);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n2584, CK => CLK, Q => 
                           REGISTERS_29_0_port, QN => n17759);
   REGISTERS_reg_30_63_inst : DFF_X1 port map( D => n2583, CK => CLK, Q => 
                           REGISTERS_30_63_port, QN => n18016);
   REGISTERS_reg_30_62_inst : DFF_X1 port map( D => n2582, CK => CLK, Q => 
                           REGISTERS_30_62_port, QN => n17080);
   REGISTERS_reg_30_61_inst : DFF_X1 port map( D => n2581, CK => CLK, Q => 
                           REGISTERS_30_61_port, QN => n17081);
   REGISTERS_reg_30_60_inst : DFF_X1 port map( D => n2580, CK => CLK, Q => 
                           REGISTERS_30_60_port, QN => n17082);
   REGISTERS_reg_30_59_inst : DFF_X1 port map( D => n2579, CK => CLK, Q => 
                           REGISTERS_30_59_port, QN => n17083);
   REGISTERS_reg_30_58_inst : DFF_X1 port map( D => n2578, CK => CLK, Q => 
                           REGISTERS_30_58_port, QN => n17159);
   REGISTERS_reg_30_57_inst : DFF_X1 port map( D => n2577, CK => CLK, Q => 
                           REGISTERS_30_57_port, QN => n17160);
   REGISTERS_reg_30_56_inst : DFF_X1 port map( D => n2576, CK => CLK, Q => 
                           REGISTERS_30_56_port, QN => n17084);
   REGISTERS_reg_30_55_inst : DFF_X1 port map( D => n2575, CK => CLK, Q => 
                           REGISTERS_30_55_port, QN => n17085);
   REGISTERS_reg_30_54_inst : DFF_X1 port map( D => n2574, CK => CLK, Q => 
                           REGISTERS_30_54_port, QN => n17086);
   REGISTERS_reg_30_53_inst : DFF_X1 port map( D => n2573, CK => CLK, Q => 
                           REGISTERS_30_53_port, QN => n17087);
   REGISTERS_reg_30_52_inst : DFF_X1 port map( D => n2572, CK => CLK, Q => 
                           REGISTERS_30_52_port, QN => n16954);
   REGISTERS_reg_30_51_inst : DFF_X1 port map( D => n2571, CK => CLK, Q => 
                           REGISTERS_30_51_port, QN => n17989);
   REGISTERS_reg_30_50_inst : DFF_X1 port map( D => n2570, CK => CLK, Q => 
                           REGISTERS_30_50_port, QN => n17990);
   REGISTERS_reg_30_49_inst : DFF_X1 port map( D => n2569, CK => CLK, Q => 
                           REGISTERS_30_49_port, QN => n17991);
   REGISTERS_reg_30_48_inst : DFF_X1 port map( D => n2568, CK => CLK, Q => 
                           REGISTERS_30_48_port, QN => n17760);
   REGISTERS_reg_30_47_inst : DFF_X1 port map( D => n2567, CK => CLK, Q => 
                           REGISTERS_30_47_port, QN => n17364);
   REGISTERS_reg_30_46_inst : DFF_X1 port map( D => n2566, CK => CLK, Q => 
                           REGISTERS_30_46_port, QN => n17365);
   REGISTERS_reg_30_45_inst : DFF_X1 port map( D => n2565, CK => CLK, Q => 
                           REGISTERS_30_45_port, QN => n17761);
   REGISTERS_reg_30_44_inst : DFF_X1 port map( D => n2564, CK => CLK, Q => 
                           REGISTERS_30_44_port, QN => n17762);
   REGISTERS_reg_30_43_inst : DFF_X1 port map( D => n2563, CK => CLK, Q => 
                           REGISTERS_30_43_port, QN => n17763);
   REGISTERS_reg_30_42_inst : DFF_X1 port map( D => n2562, CK => CLK, Q => 
                           REGISTERS_30_42_port, QN => n17992);
   REGISTERS_reg_30_41_inst : DFF_X1 port map( D => n2561, CK => CLK, Q => 
                           REGISTERS_30_41_port, QN => n17993);
   REGISTERS_reg_30_40_inst : DFF_X1 port map( D => n2560, CK => CLK, Q => 
                           REGISTERS_30_40_port, QN => n17994);
   REGISTERS_reg_30_39_inst : DFF_X1 port map( D => n2559, CK => CLK, Q => 
                           REGISTERS_30_39_port, QN => n17995);
   REGISTERS_reg_30_38_inst : DFF_X1 port map( D => n2558, CK => CLK, Q => 
                           REGISTERS_30_38_port, QN => n17996);
   REGISTERS_reg_30_37_inst : DFF_X1 port map( D => n2557, CK => CLK, Q => 
                           REGISTERS_30_37_port, QN => n17366);
   REGISTERS_reg_30_36_inst : DFF_X1 port map( D => n2556, CK => CLK, Q => 
                           REGISTERS_30_36_port, QN => n17764);
   REGISTERS_reg_30_35_inst : DFF_X1 port map( D => n2555, CK => CLK, Q => 
                           REGISTERS_30_35_port, QN => n17997);
   REGISTERS_reg_30_34_inst : DFF_X1 port map( D => n2554, CK => CLK, Q => 
                           REGISTERS_30_34_port, QN => n17998);
   REGISTERS_reg_30_33_inst : DFF_X1 port map( D => n2553, CK => CLK, Q => 
                           REGISTERS_30_33_port, QN => n17367);
   REGISTERS_reg_30_32_inst : DFF_X1 port map( D => n2552, CK => CLK, Q => 
                           REGISTERS_30_32_port, QN => n17368);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n2551, CK => CLK, Q => 
                           REGISTERS_30_31_port, QN => n17369);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n2550, CK => CLK, Q => 
                           REGISTERS_30_30_port, QN => n17999);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n2549, CK => CLK, Q => 
                           REGISTERS_30_29_port, QN => n18000);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n2548, CK => CLK, Q => 
                           REGISTERS_30_28_port, QN => n17765);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n2547, CK => CLK, Q => 
                           REGISTERS_30_27_port, QN => n17088);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n2546, CK => CLK, Q => 
                           REGISTERS_30_26_port, QN => n16955);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n2545, CK => CLK, Q => 
                           REGISTERS_30_25_port, QN => n17161);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n2544, CK => CLK, Q => 
                           REGISTERS_30_24_port, QN => n17089);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n2543, CK => CLK, Q => 
                           REGISTERS_30_23_port, QN => n17162);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n2542, CK => CLK, Q => 
                           REGISTERS_30_22_port, QN => n16956);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n2541, CK => CLK, Q => 
                           REGISTERS_30_21_port, QN => n17090);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n2540, CK => n13730, Q => 
                           REGISTERS_30_20_port, QN => n17163);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n2539, CK => CLK, Q => 
                           REGISTERS_30_19_port, QN => n17091);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n2538, CK => CLK, Q => 
                           REGISTERS_30_18_port, QN => n16957);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n2537, CK => CLK, Q => 
                           REGISTERS_30_17_port, QN => n17092);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n2536, CK => CLK, Q => 
                           REGISTERS_30_16_port, QN => n17164);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n2535, CK => CLK, Q => 
                           REGISTERS_30_15_port, QN => n17370);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n2534, CK => CLK, Q => 
                           REGISTERS_30_14_port, QN => n17766);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n2533, CK => CLK, Q => 
                           REGISTERS_30_13_port, QN => n17371);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n2532, CK => CLK, Q => 
                           REGISTERS_30_12_port, QN => n17767);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n2531, CK => CLK, Q => 
                           REGISTERS_30_11_port, QN => n17768);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n2530, CK => CLK, Q => 
                           REGISTERS_30_10_port, QN => n17372);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n2529, CK => CLK, Q => 
                           REGISTERS_30_9_port, QN => n17769);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n2528, CK => CLK, Q => 
                           REGISTERS_30_8_port, QN => n17770);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n2527, CK => CLK, Q => 
                           REGISTERS_30_7_port, QN => n17771);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n2526, CK => CLK, Q => 
                           REGISTERS_30_6_port, QN => n17772);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n2525, CK => CLK, Q => 
                           REGISTERS_30_5_port, QN => n18001);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n2524, CK => CLK, Q => 
                           REGISTERS_30_4_port, QN => n17773);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n2523, CK => CLK, Q => 
                           REGISTERS_30_3_port, QN => n17774);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n2522, CK => CLK, Q => 
                           REGISTERS_30_2_port, QN => n17373);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n2521, CK => CLK, Q => 
                           REGISTERS_30_1_port, QN => n17775);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n2520, CK => CLK, Q => 
                           REGISTERS_30_0_port, QN => n17776);
   REGISTERS_reg_31_63_inst : DFF_X1 port map( D => n2519, CK => CLK, Q => 
                           REGISTERS_31_63_port, QN => n18242);
   REGISTERS_reg_31_62_inst : DFF_X1 port map( D => n2518, CK => CLK, Q => 
                           REGISTERS_31_62_port, QN => n17093);
   REGISTERS_reg_31_61_inst : DFF_X1 port map( D => n2517, CK => CLK, Q => 
                           REGISTERS_31_61_port, QN => n17094);
   REGISTERS_reg_31_60_inst : DFF_X1 port map( D => n2516, CK => CLK, Q => 
                           REGISTERS_31_60_port, QN => n16958);
   REGISTERS_reg_31_59_inst : DFF_X1 port map( D => n2515, CK => CLK, Q => 
                           REGISTERS_31_59_port, QN => n17165);
   REGISTERS_reg_31_58_inst : DFF_X1 port map( D => n2514, CK => CLK, Q => 
                           REGISTERS_31_58_port, QN => n17095);
   REGISTERS_reg_31_57_inst : DFF_X1 port map( D => n2513, CK => CLK, Q => 
                           REGISTERS_31_57_port, QN => n16959);
   REGISTERS_reg_31_56_inst : DFF_X1 port map( D => n2512, CK => CLK, Q => 
                           REGISTERS_31_56_port, QN => n17166);
   REGISTERS_reg_31_55_inst : DFF_X1 port map( D => n2511, CK => CLK, Q => 
                           REGISTERS_31_55_port, QN => n17167);
   REGISTERS_reg_31_54_inst : DFF_X1 port map( D => n2510, CK => CLK, Q => 
                           REGISTERS_31_54_port, QN => n17096);
   REGISTERS_reg_31_53_inst : DFF_X1 port map( D => n2509, CK => CLK, Q => 
                           REGISTERS_31_53_port, QN => n16960);
   REGISTERS_reg_31_52_inst : DFF_X1 port map( D => n2508, CK => CLK, Q => 
                           REGISTERS_31_52_port, QN => n17097);
   REGISTERS_reg_31_51_inst : DFF_X1 port map( D => n2507, CK => CLK, Q => 
                           REGISTERS_31_51_port, QN => n17777);
   REGISTERS_reg_31_50_inst : DFF_X1 port map( D => n2506, CK => CLK, Q => 
                           REGISTERS_31_50_port, QN => n17778);
   REGISTERS_reg_31_49_inst : DFF_X1 port map( D => n2505, CK => CLK, Q => 
                           REGISTERS_31_49_port, QN => n17779);
   REGISTERS_reg_31_48_inst : DFF_X1 port map( D => n2504, CK => n13730, Q => 
                           REGISTERS_31_48_port, QN => n18002);
   REGISTERS_reg_31_47_inst : DFF_X1 port map( D => n2503, CK => CLK, Q => 
                           REGISTERS_31_47_port, QN => n17374);
   REGISTERS_reg_31_46_inst : DFF_X1 port map( D => n2502, CK => CLK, Q => 
                           REGISTERS_31_46_port, QN => n17375);
   REGISTERS_reg_31_45_inst : DFF_X1 port map( D => n2501, CK => CLK, Q => 
                           REGISTERS_31_45_port, QN => n17376);
   REGISTERS_reg_31_44_inst : DFF_X1 port map( D => n2500, CK => CLK, Q => 
                           REGISTERS_31_44_port, QN => n17377);
   REGISTERS_reg_31_43_inst : DFF_X1 port map( D => n2499, CK => CLK, Q => 
                           REGISTERS_31_43_port, QN => n17378);
   REGISTERS_reg_31_42_inst : DFF_X1 port map( D => n2498, CK => CLK, Q => 
                           REGISTERS_31_42_port, QN => n17780);
   REGISTERS_reg_31_41_inst : DFF_X1 port map( D => n2497, CK => CLK, Q => 
                           REGISTERS_31_41_port, QN => n17379);
   REGISTERS_reg_31_40_inst : DFF_X1 port map( D => n2496, CK => CLK, Q => 
                           REGISTERS_31_40_port, QN => n18003);
   REGISTERS_reg_31_39_inst : DFF_X1 port map( D => n2495, CK => CLK, Q => 
                           REGISTERS_31_39_port, QN => n17781);
   REGISTERS_reg_31_38_inst : DFF_X1 port map( D => n2494, CK => CLK, Q => 
                           REGISTERS_31_38_port, QN => n17782);
   REGISTERS_reg_31_37_inst : DFF_X1 port map( D => n2493, CK => CLK, Q => 
                           REGISTERS_31_37_port, QN => n17380);
   REGISTERS_reg_31_36_inst : DFF_X1 port map( D => n2492, CK => CLK, Q => 
                           REGISTERS_31_36_port, QN => n17783);
   REGISTERS_reg_31_35_inst : DFF_X1 port map( D => n2491, CK => CLK, Q => 
                           REGISTERS_31_35_port, QN => n17784);
   REGISTERS_reg_31_34_inst : DFF_X1 port map( D => n2490, CK => CLK, Q => 
                           REGISTERS_31_34_port, QN => n17381);
   REGISTERS_reg_31_33_inst : DFF_X1 port map( D => n2489, CK => CLK, Q => 
                           REGISTERS_31_33_port, QN => n17382);
   REGISTERS_reg_31_32_inst : DFF_X1 port map( D => n2488, CK => CLK, Q => 
                           REGISTERS_31_32_port, QN => n17383);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n2487, CK => CLK, Q => 
                           REGISTERS_31_31_port, QN => n17384);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n2486, CK => CLK, Q => 
                           REGISTERS_31_30_port, QN => n17385);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n2485, CK => CLK, Q => 
                           REGISTERS_31_29_port, QN => n17785);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n2484, CK => CLK, Q => 
                           REGISTERS_31_28_port, QN => n17786);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n2483, CK => CLK, Q => 
                           REGISTERS_31_27_port, QN => n17098);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n2482, CK => CLK, Q => 
                           REGISTERS_31_26_port, QN => n17099);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n2481, CK => CLK, Q => 
                           REGISTERS_31_25_port, QN => n16961);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n2480, CK => CLK, Q => 
                           REGISTERS_31_24_port, QN => n17168);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n2479, CK => CLK, Q => 
                           REGISTERS_31_23_port, QN => n17100);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n2478, CK => CLK, Q => 
                           REGISTERS_31_22_port, QN => n17101);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n2477, CK => CLK, Q => 
                           REGISTERS_31_21_port, QN => n17102);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n2476, CK => CLK, Q => 
                           REGISTERS_31_20_port, QN => n17103);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n2475, CK => CLK, Q => 
                           REGISTERS_31_19_port, QN => n16962);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n2474, CK => CLK, Q => 
                           REGISTERS_31_18_port, QN => n17169);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n2473, CK => CLK, Q => 
                           REGISTERS_31_17_port, QN => n17104);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n2472, CK => CLK, Q => 
                           REGISTERS_31_16_port, QN => n17170);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n2471, CK => CLK, Q => 
                           REGISTERS_31_15_port, QN => n17787);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n2470, CK => CLK, Q => 
                           REGISTERS_31_14_port, QN => n17386);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n2469, CK => CLK, Q => 
                           REGISTERS_31_13_port, QN => n17788);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n2468, CK => CLK, Q => 
                           REGISTERS_31_12_port, QN => n18004);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n2467, CK => CLK, Q => 
                           REGISTERS_31_11_port, QN => n18005);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n2466, CK => CLK, Q => 
                           REGISTERS_31_10_port, QN => n18006);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n2465, CK => CLK, Q => 
                           REGISTERS_31_9_port, QN => n18007);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n2464, CK => CLK, Q => 
                           REGISTERS_31_8_port, QN => n17789);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n2463, CK => CLK, Q => 
                           REGISTERS_31_7_port, QN => n18008);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n2462, CK => CLK, Q => 
                           REGISTERS_31_6_port, QN => n17387);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n2461, CK => CLK, Q => 
                           REGISTERS_31_5_port, QN => n17790);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n2460, CK => CLK, Q => 
                           REGISTERS_31_4_port, QN => n18009);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n2459, CK => CLK, Q => 
                           REGISTERS_31_3_port, QN => n18010);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n2458, CK => CLK, Q => 
                           REGISTERS_31_2_port, QN => n17791);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n2457, CK => CLK, Q => 
                           REGISTERS_31_1_port, QN => n17792);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n2456, CK => CLK, Q => 
                           REGISTERS_31_0_port, QN => n17793);
   out1_signal_reg_63_inst : DFF_X1 port map( D => n8506, CK => CLK, Q => 
                           OUT1(63), QN => n8505);
   out1_signal_reg_62_inst : DFF_X1 port map( D => n8507, CK => CLK, Q => 
                           OUT1(62), QN => n8504);
   out1_signal_reg_61_inst : DFF_X1 port map( D => n8508, CK => CLK, Q => 
                           OUT1(61), QN => n8503);
   out1_signal_reg_60_inst : DFF_X1 port map( D => n8509, CK => CLK, Q => 
                           OUT1(60), QN => n8502);
   out1_signal_reg_59_inst : DFF_X1 port map( D => n8510, CK => CLK, Q => 
                           OUT1(59), QN => n8501);
   out1_signal_reg_58_inst : DFF_X1 port map( D => n8511, CK => CLK, Q => 
                           OUT1(58), QN => n8500);
   out1_signal_reg_57_inst : DFF_X1 port map( D => n8512, CK => CLK, Q => 
                           OUT1(57), QN => n8499);
   out1_signal_reg_56_inst : DFF_X1 port map( D => n8513, CK => CLK, Q => 
                           OUT1(56), QN => n8498);
   out1_signal_reg_55_inst : DFF_X1 port map( D => n8514, CK => CLK, Q => 
                           OUT1(55), QN => n8497);
   out1_signal_reg_54_inst : DFF_X1 port map( D => n8515, CK => CLK, Q => 
                           OUT1(54), QN => n8496);
   out1_signal_reg_53_inst : DFF_X1 port map( D => n8516, CK => CLK, Q => 
                           OUT1(53), QN => n8495);
   out1_signal_reg_52_inst : DFF_X1 port map( D => n8517, CK => CLK, Q => 
                           OUT1(52), QN => n8494);
   out1_signal_reg_51_inst : DFF_X1 port map( D => n8518, CK => CLK, Q => 
                           OUT1(51), QN => n8493);
   out1_signal_reg_50_inst : DFF_X1 port map( D => n8519, CK => CLK, Q => 
                           OUT1(50), QN => n8492);
   out1_signal_reg_49_inst : DFF_X1 port map( D => n8520, CK => CLK, Q => 
                           OUT1(49), QN => n8491);
   out1_signal_reg_48_inst : DFF_X1 port map( D => n8521, CK => CLK, Q => 
                           OUT1(48), QN => n8490);
   out1_signal_reg_47_inst : DFF_X1 port map( D => n8522, CK => CLK, Q => 
                           OUT1(47), QN => n8489);
   out1_signal_reg_46_inst : DFF_X1 port map( D => n8523, CK => CLK, Q => 
                           OUT1(46), QN => n8488);
   out1_signal_reg_45_inst : DFF_X1 port map( D => n8524, CK => CLK, Q => 
                           OUT1(45), QN => n8487);
   out1_signal_reg_44_inst : DFF_X1 port map( D => n8525, CK => CLK, Q => 
                           OUT1(44), QN => n8486);
   out1_signal_reg_43_inst : DFF_X1 port map( D => n8526, CK => CLK, Q => 
                           OUT1(43), QN => n8485);
   out1_signal_reg_42_inst : DFF_X1 port map( D => n8527, CK => CLK, Q => 
                           OUT1(42), QN => n8484);
   out1_signal_reg_41_inst : DFF_X1 port map( D => n8528, CK => CLK, Q => 
                           OUT1(41), QN => n8483);
   out1_signal_reg_40_inst : DFF_X1 port map( D => n8529, CK => CLK, Q => 
                           OUT1(40), QN => n8482);
   out1_signal_reg_39_inst : DFF_X1 port map( D => n8530, CK => CLK, Q => 
                           OUT1(39), QN => n8481);
   out1_signal_reg_38_inst : DFF_X1 port map( D => n8531, CK => CLK, Q => 
                           OUT1(38), QN => n8480);
   out1_signal_reg_37_inst : DFF_X1 port map( D => n8532, CK => CLK, Q => 
                           OUT1(37), QN => n8479);
   out1_signal_reg_36_inst : DFF_X1 port map( D => n8533, CK => CLK, Q => 
                           OUT1(36), QN => n8478);
   out1_signal_reg_35_inst : DFF_X1 port map( D => n8534, CK => CLK, Q => 
                           OUT1(35), QN => n8477);
   out1_signal_reg_34_inst : DFF_X1 port map( D => n8535, CK => CLK, Q => 
                           OUT1(34), QN => n8476);
   out1_signal_reg_33_inst : DFF_X1 port map( D => n8536, CK => CLK, Q => 
                           OUT1(33), QN => n8475);
   out1_signal_reg_32_inst : DFF_X1 port map( D => n8537, CK => CLK, Q => 
                           OUT1(32), QN => n8474);
   out1_signal_reg_31_inst : DFF_X1 port map( D => n8538, CK => CLK, Q => 
                           OUT1(31), QN => n8473);
   out1_signal_reg_30_inst : DFF_X1 port map( D => n8539, CK => CLK, Q => 
                           OUT1(30), QN => n8472);
   out1_signal_reg_29_inst : DFF_X1 port map( D => n8540, CK => CLK, Q => 
                           OUT1(29), QN => n8471);
   out1_signal_reg_28_inst : DFF_X1 port map( D => n8541, CK => CLK, Q => 
                           OUT1(28), QN => n8470);
   out1_signal_reg_27_inst : DFF_X1 port map( D => n8542, CK => CLK, Q => 
                           OUT1(27), QN => n8469);
   out1_signal_reg_26_inst : DFF_X1 port map( D => n8543, CK => CLK, Q => 
                           OUT1(26), QN => n8468);
   out1_signal_reg_25_inst : DFF_X1 port map( D => n8544, CK => CLK, Q => 
                           OUT1(25), QN => n8467);
   out1_signal_reg_24_inst : DFF_X1 port map( D => n8545, CK => CLK, Q => 
                           OUT1(24), QN => n8466);
   out1_signal_reg_23_inst : DFF_X1 port map( D => n8546, CK => CLK, Q => 
                           OUT1(23), QN => n8465);
   out1_signal_reg_22_inst : DFF_X1 port map( D => n8547, CK => CLK, Q => 
                           OUT1(22), QN => n8464);
   out1_signal_reg_21_inst : DFF_X1 port map( D => n8548, CK => CLK, Q => 
                           OUT1(21), QN => n8463);
   out1_signal_reg_20_inst : DFF_X1 port map( D => n8549, CK => CLK, Q => 
                           OUT1(20), QN => n8462);
   out1_signal_reg_19_inst : DFF_X1 port map( D => n8550, CK => CLK, Q => 
                           OUT1(19), QN => n8461);
   out1_signal_reg_18_inst : DFF_X1 port map( D => n8551, CK => CLK, Q => 
                           OUT1(18), QN => n8460);
   out1_signal_reg_17_inst : DFF_X1 port map( D => n8552, CK => CLK, Q => 
                           OUT1(17), QN => n8459);
   out1_signal_reg_16_inst : DFF_X1 port map( D => n8553, CK => CLK, Q => 
                           OUT1(16), QN => n8458);
   out1_signal_reg_15_inst : DFF_X1 port map( D => n8554, CK => CLK, Q => 
                           OUT1(15), QN => n8457);
   out1_signal_reg_14_inst : DFF_X1 port map( D => n8555, CK => CLK, Q => 
                           OUT1(14), QN => n8456);
   out1_signal_reg_13_inst : DFF_X1 port map( D => n8556, CK => CLK, Q => 
                           OUT1(13), QN => n8455);
   out1_signal_reg_12_inst : DFF_X1 port map( D => n8557, CK => CLK, Q => 
                           OUT1(12), QN => n8454);
   out1_signal_reg_11_inst : DFF_X1 port map( D => n8558, CK => CLK, Q => 
                           OUT1(11), QN => n8453);
   out1_signal_reg_10_inst : DFF_X1 port map( D => n8559, CK => CLK, Q => 
                           OUT1(10), QN => n8452);
   out1_signal_reg_9_inst : DFF_X1 port map( D => n8560, CK => CLK, Q => 
                           OUT1(9), QN => n8451);
   out1_signal_reg_8_inst : DFF_X1 port map( D => n8561, CK => CLK, Q => 
                           OUT1(8), QN => n8450);
   out1_signal_reg_7_inst : DFF_X1 port map( D => n8562, CK => CLK, Q => 
                           OUT1(7), QN => n8449);
   out1_signal_reg_6_inst : DFF_X1 port map( D => n8563, CK => CLK, Q => 
                           OUT1(6), QN => n8448);
   out1_signal_reg_5_inst : DFF_X1 port map( D => n8564, CK => CLK, Q => 
                           OUT1(5), QN => n8447);
   out1_signal_reg_4_inst : DFF_X1 port map( D => n8565, CK => CLK, Q => 
                           OUT1(4), QN => n8446);
   out1_signal_reg_3_inst : DFF_X1 port map( D => n8566, CK => CLK, Q => 
                           OUT1(3), QN => n8445);
   out1_signal_reg_2_inst : DFF_X1 port map( D => n8567, CK => CLK, Q => 
                           OUT1(2), QN => n8444);
   out1_signal_reg_1_inst : DFF_X1 port map( D => n8568, CK => CLK, Q => 
                           OUT1(1), QN => n8443);
   out1_signal_reg_0_inst : DFF_X1 port map( D => n8569, CK => CLK, Q => 
                           OUT1(0), QN => n8442);
   out2_signal_reg_63_inst : DFF_X1 port map( D => n8570, CK => CLK, Q => 
                           OUT2(63), QN => n8441);
   out2_signal_reg_62_inst : DFF_X1 port map( D => n8571, CK => CLK, Q => 
                           OUT2(62), QN => n8440);
   out2_signal_reg_61_inst : DFF_X1 port map( D => n8572, CK => CLK, Q => 
                           OUT2(61), QN => n8439);
   out2_signal_reg_60_inst : DFF_X1 port map( D => n8573, CK => CLK, Q => 
                           OUT2(60), QN => n8438);
   out2_signal_reg_59_inst : DFF_X1 port map( D => n8574, CK => CLK, Q => 
                           OUT2(59), QN => n8437);
   out2_signal_reg_58_inst : DFF_X1 port map( D => n8575, CK => CLK, Q => 
                           OUT2(58), QN => n8436);
   out2_signal_reg_57_inst : DFF_X1 port map( D => n8576, CK => CLK, Q => 
                           OUT2(57), QN => n8435);
   out2_signal_reg_56_inst : DFF_X1 port map( D => n8577, CK => CLK, Q => 
                           OUT2(56), QN => n8434);
   out2_signal_reg_55_inst : DFF_X1 port map( D => n8578, CK => CLK, Q => 
                           OUT2(55), QN => n8433);
   out2_signal_reg_54_inst : DFF_X1 port map( D => n8579, CK => CLK, Q => 
                           OUT2(54), QN => n8432);
   out2_signal_reg_53_inst : DFF_X1 port map( D => n8580, CK => CLK, Q => 
                           OUT2(53), QN => n8431);
   out2_signal_reg_52_inst : DFF_X1 port map( D => n8581, CK => CLK, Q => 
                           OUT2(52), QN => n8430);
   out2_signal_reg_51_inst : DFF_X1 port map( D => n8582, CK => CLK, Q => 
                           OUT2(51), QN => n8429);
   out2_signal_reg_50_inst : DFF_X1 port map( D => n8583, CK => CLK, Q => 
                           OUT2(50), QN => n8428);
   out2_signal_reg_49_inst : DFF_X1 port map( D => n8584, CK => CLK, Q => 
                           OUT2(49), QN => n8427);
   out2_signal_reg_48_inst : DFF_X1 port map( D => n8585, CK => CLK, Q => 
                           OUT2(48), QN => n8426);
   out2_signal_reg_47_inst : DFF_X1 port map( D => n8586, CK => CLK, Q => 
                           OUT2(47), QN => n8425);
   out2_signal_reg_46_inst : DFF_X1 port map( D => n8587, CK => CLK, Q => 
                           OUT2(46), QN => n8424);
   out2_signal_reg_45_inst : DFF_X1 port map( D => n8588, CK => CLK, Q => 
                           OUT2(45), QN => n8423);
   out2_signal_reg_44_inst : DFF_X1 port map( D => n8589, CK => CLK, Q => 
                           OUT2(44), QN => n8422);
   out2_signal_reg_43_inst : DFF_X1 port map( D => n8590, CK => CLK, Q => 
                           OUT2(43), QN => n8421);
   out2_signal_reg_42_inst : DFF_X1 port map( D => n8591, CK => CLK, Q => 
                           OUT2(42), QN => n8420);
   out2_signal_reg_41_inst : DFF_X1 port map( D => n8592, CK => CLK, Q => 
                           OUT2(41), QN => n8419);
   out2_signal_reg_40_inst : DFF_X1 port map( D => n8593, CK => CLK, Q => 
                           OUT2(40), QN => n8418);
   out2_signal_reg_39_inst : DFF_X1 port map( D => n8594, CK => CLK, Q => 
                           OUT2(39), QN => n8417);
   out2_signal_reg_38_inst : DFF_X1 port map( D => n8595, CK => CLK, Q => 
                           OUT2(38), QN => n8416);
   out2_signal_reg_37_inst : DFF_X1 port map( D => n8596, CK => CLK, Q => 
                           OUT2(37), QN => n8415);
   out2_signal_reg_36_inst : DFF_X1 port map( D => n8597, CK => CLK, Q => 
                           OUT2(36), QN => n8414);
   out2_signal_reg_35_inst : DFF_X1 port map( D => n8598, CK => CLK, Q => 
                           OUT2(35), QN => n8413);
   out2_signal_reg_34_inst : DFF_X1 port map( D => n8599, CK => CLK, Q => 
                           OUT2(34), QN => n8412);
   out2_signal_reg_33_inst : DFF_X1 port map( D => n8600, CK => CLK, Q => 
                           OUT2(33), QN => n8411);
   out2_signal_reg_32_inst : DFF_X1 port map( D => n8601, CK => CLK, Q => 
                           OUT2(32), QN => n8410);
   out2_signal_reg_31_inst : DFF_X1 port map( D => n8602, CK => CLK, Q => 
                           OUT2(31), QN => n8409);
   out2_signal_reg_30_inst : DFF_X1 port map( D => n8603, CK => CLK, Q => 
                           OUT2(30), QN => n8408);
   out2_signal_reg_29_inst : DFF_X1 port map( D => n8604, CK => CLK, Q => 
                           OUT2(29), QN => n8407);
   out2_signal_reg_28_inst : DFF_X1 port map( D => n8605, CK => CLK, Q => 
                           OUT2(28), QN => n8406);
   out2_signal_reg_27_inst : DFF_X1 port map( D => n8606, CK => CLK, Q => 
                           OUT2(27), QN => n8405);
   out2_signal_reg_26_inst : DFF_X1 port map( D => n8607, CK => CLK, Q => 
                           OUT2(26), QN => n8404);
   out2_signal_reg_25_inst : DFF_X1 port map( D => n8608, CK => CLK, Q => 
                           OUT2(25), QN => n8403);
   out2_signal_reg_24_inst : DFF_X1 port map( D => n8609, CK => CLK, Q => 
                           OUT2(24), QN => n8402);
   out2_signal_reg_23_inst : DFF_X1 port map( D => n8610, CK => CLK, Q => 
                           OUT2(23), QN => n8401);
   out2_signal_reg_22_inst : DFF_X1 port map( D => n8611, CK => CLK, Q => 
                           OUT2(22), QN => n8400);
   out2_signal_reg_21_inst : DFF_X1 port map( D => n8612, CK => CLK, Q => 
                           OUT2(21), QN => n8399);
   out2_signal_reg_20_inst : DFF_X1 port map( D => n8613, CK => CLK, Q => 
                           OUT2(20), QN => n8398);
   out2_signal_reg_19_inst : DFF_X1 port map( D => n8614, CK => CLK, Q => 
                           OUT2(19), QN => n8397);
   out2_signal_reg_18_inst : DFF_X1 port map( D => n8615, CK => CLK, Q => 
                           OUT2(18), QN => n8396);
   out2_signal_reg_17_inst : DFF_X1 port map( D => n8616, CK => CLK, Q => 
                           OUT2(17), QN => n8395);
   out2_signal_reg_16_inst : DFF_X1 port map( D => n8617, CK => CLK, Q => 
                           OUT2(16), QN => n8394);
   out2_signal_reg_15_inst : DFF_X1 port map( D => n8618, CK => CLK, Q => 
                           OUT2(15), QN => n8393);
   out2_signal_reg_14_inst : DFF_X1 port map( D => n8619, CK => CLK, Q => 
                           OUT2(14), QN => n8392);
   out2_signal_reg_13_inst : DFF_X1 port map( D => n8620, CK => CLK, Q => 
                           OUT2(13), QN => n8391);
   out2_signal_reg_12_inst : DFF_X1 port map( D => n8621, CK => CLK, Q => 
                           OUT2(12), QN => n8390);
   out2_signal_reg_11_inst : DFF_X1 port map( D => n8622, CK => CLK, Q => 
                           OUT2(11), QN => n8389);
   out2_signal_reg_10_inst : DFF_X1 port map( D => n8623, CK => CLK, Q => 
                           OUT2(10), QN => n8388);
   out2_signal_reg_9_inst : DFF_X1 port map( D => n8624, CK => CLK, Q => 
                           OUT2(9), QN => n8387);
   out2_signal_reg_8_inst : DFF_X1 port map( D => n8625, CK => CLK, Q => 
                           OUT2(8), QN => n8386);
   out2_signal_reg_7_inst : DFF_X1 port map( D => n8626, CK => CLK, Q => 
                           OUT2(7), QN => n8385);
   out2_signal_reg_6_inst : DFF_X1 port map( D => n8627, CK => CLK, Q => 
                           OUT2(6), QN => n8384);
   out2_signal_reg_5_inst : DFF_X1 port map( D => n8628, CK => CLK, Q => 
                           OUT2(5), QN => n8383);
   out2_signal_reg_4_inst : DFF_X1 port map( D => n8629, CK => CLK, Q => 
                           OUT2(4), QN => n8382);
   out2_signal_reg_3_inst : DFF_X1 port map( D => n8630, CK => CLK, Q => 
                           OUT2(3), QN => n8381);
   out2_signal_reg_2_inst : DFF_X1 port map( D => n8631, CK => CLK, Q => 
                           OUT2(2), QN => n8380);
   out2_signal_reg_1_inst : DFF_X1 port map( D => n8632, CK => CLK, Q => 
                           OUT2(1), QN => n8379);
   out2_signal_reg_0_inst : DFF_X1 port map( D => n8633, CK => CLK, Q => 
                           OUT2(0), QN => n8378);
   U11778 : CLKBUF_X1 port map( A => CLK, Z => n13730);
   U11779 : NOR3_X2 port map( A1 => ADD_WR(3), A2 => n16678, A3 => n16644, ZN 
                           => n16639);
   U11780 : INV_X8 port map( A => RESET, ZN => n13731);
   U11781 : BUF_X4 port map( A => n13761, Z => n15154);
   U11782 : BUF_X4 port map( A => n13760, Z => n15128);
   U11783 : BUF_X4 port map( A => n13758, Z => n15144);
   U11784 : BUF_X4 port map( A => n13754, Z => n15142);
   U11785 : BUF_X4 port map( A => n13759, Z => n15126);
   U11786 : BUF_X4 port map( A => n13757, Z => n15145);
   U11787 : BUF_X4 port map( A => n13755, Z => n15150);
   U11788 : BUF_X4 port map( A => n13748, Z => n15152);
   U11789 : BUF_X4 port map( A => n13747, Z => n15130);
   U11790 : BUF_X4 port map( A => n13746, Z => n15127);
   U11791 : BUF_X4 port map( A => n13743, Z => n15156);
   U11792 : BUF_X4 port map( A => n13745, Z => n15132);
   U11793 : BUF_X4 port map( A => n13741, Z => n15140);
   U11794 : BUF_X4 port map( A => n13744, Z => n15153);
   U11795 : BUF_X4 port map( A => n13740, Z => n15138);
   U11796 : BUF_X4 port map( A => n15183, Z => n16574);
   U11797 : BUF_X4 port map( A => n15171, Z => n16555);
   U11798 : BUF_X4 port map( A => n15197, Z => n16569);
   U11799 : BUF_X4 port map( A => n15203, Z => n16561);
   U11800 : BUF_X4 port map( A => n15174, Z => n16580);
   U11801 : BUF_X4 port map( A => n15169, Z => n16581);
   U11802 : BUF_X4 port map( A => n15196, Z => n16556);
   U11803 : BUF_X4 port map( A => n15170, Z => n16557);
   U11804 : BUF_X4 port map( A => n15198, Z => n16573);
   U11805 : BUF_X4 port map( A => n15173, Z => n16560);
   U11806 : BUF_X4 port map( A => n15205, Z => n16571);
   U11807 : BUF_X4 port map( A => n15182, Z => n16570);
   U11808 : BUF_X4 port map( A => n15187, Z => n16558);
   U11809 : BUF_X4 port map( A => n15200, Z => n16583);
   U11810 : BUF_X4 port map( A => n15172, Z => n16579);
   U11811 : BUF_X4 port map( A => n15181, Z => n16562);
   U11812 : BUF_X4 port map( A => n15186, Z => n16572);
   U11813 : BUF_X4 port map( A => n15195, Z => n16584);
   U11814 : BUF_X4 port map( A => n15180, Z => n16582);
   U11815 : BUF_X4 port map( A => n15190, Z => n16559);
   U11816 : BUF_X4 port map( A => n13775, Z => n15143);
   U11817 : BUF_X4 port map( A => n15201, Z => n16567);
   U11818 : BUF_X4 port map( A => n15175, Z => n16568);
   U11819 : BUF_X4 port map( A => n13767, Z => n15157);
   U11820 : BUF_X4 port map( A => n13769, Z => n15129);
   U11821 : NOR3_X2 port map( A1 => ADD_WR(3), A2 => n16678, A3 => n16712, ZN 
                           => n16707);
   U11822 : INV_X1 port map( A => n13770, ZN => n14506);
   U11823 : INV_X1 port map( A => n16216, ZN => n15366);
   U11824 : INV_X1 port map( A => n16344, ZN => n15258);
   U11825 : INV_X1 port map( A => n16215, ZN => n15344);
   U11826 : OR3_X1 port map( A1 => n15184, A2 => ADD_RD2(1), A3 => ADD_RD2(0), 
                           ZN => n15236);
   U11827 : CLKBUF_X1 port map( A => n14910, Z => n16049);
   U11828 : INV_X1 port map( A => n16322, ZN => n15556);
   U11829 : INV_X1 port map( A => n15746, ZN => n15301);
   U11830 : OR2_X1 port map( A1 => n13735, A2 => n13732, ZN => n14461);
   U11831 : OR2_X1 port map( A1 => ADD_RD1(1), A2 => n13732, ZN => n13785);
   U11832 : INV_X1 port map( A => ADD_RD2(4), ZN => n15168);
   U11833 : OR2_X1 port map( A1 => n13742, A2 => ADD_RD1(3), ZN => n13772);
   U11834 : INV_X1 port map( A => ADD_RD1(0), ZN => n13734);
   U11835 : INV_X1 port map( A => ADD_RD2(2), ZN => n15184);
   U11836 : CLKBUF_X1 port map( A => n14837, Z => n15096);
   U11837 : INV_X1 port map( A => n15556, ZN => n16430);
   U11838 : INV_X1 port map( A => n15366, ZN => n16594);
   U11839 : CLKBUF_X1 port map( A => n16545, Z => n16596);
   U11840 : INV_X1 port map( A => n15344, ZN => n16542);
   U11841 : CLKBUF_X1 port map( A => n16547, Z => n16597);
   U11842 : INV_X1 port map( A => n15301, ZN => n16593);
   U11843 : INV_X1 port map( A => n15258, ZN => n16592);
   U11844 : CLKBUF_X1 port map( A => n15089, Z => n15116);
   U11845 : INV_X1 port map( A => n14461, ZN => n15119);
   U11846 : CLKBUF_X1 port map( A => n14506, Z => n15019);
   U11847 : INV_X1 port map( A => n13785, ZN => n15118);
   U11848 : CLKBUF_X1 port map( A => n14506, Z => n14759);
   U11849 : CLKBUF_X1 port map( A => n15065, Z => n15120);
   U11850 : INV_X1 port map( A => n13773, ZN => n15090);
   U11851 : CLKBUF_X1 port map( A => n15043, Z => n14781);
   U11852 : INV_X1 port map( A => n13753, ZN => n15117);
   U11853 : INV_X1 port map( A => ENABLE, ZN => n16678);
   U11854 : AND4_X1 port map( A1 => n16601, A2 => n16600, A3 => n16599, A4 => 
                           n16598, ZN => n16602);
   U11855 : AND4_X1 port map( A1 => n16434, A2 => n16433, A3 => n16432, A4 => 
                           n16431, ZN => n16435);
   U11856 : AND4_X1 port map( A1 => n16283, A2 => n16282, A3 => n16281, A4 => 
                           n16280, ZN => n16284);
   U11857 : AND4_X1 port map( A1 => n16113, A2 => n16112, A3 => n16111, A4 => 
                           n16110, ZN => n16114);
   U11858 : CLKBUF_X1 port map( A => n16553, Z => n16603);
   U11859 : AND4_X1 port map( A1 => n15815, A2 => n15814, A3 => n15813, A4 => 
                           n15812, ZN => n15816);
   U11860 : AND4_X1 port map( A1 => n15665, A2 => n15664, A3 => n15663, A4 => 
                           n15662, ZN => n15666);
   U11861 : AND4_X1 port map( A1 => n15517, A2 => n15516, A3 => n15515, A4 => 
                           n15514, ZN => n15518);
   U11862 : AND4_X1 port map( A1 => n15348, A2 => n15347, A3 => n15346, A4 => 
                           n15345, ZN => n15349);
   U11863 : AND4_X1 port map( A1 => n15218, A2 => n15217, A3 => n15216, A4 => 
                           n15215, ZN => n15219);
   U11864 : AND4_X1 port map( A1 => n15000, A2 => n14999, A3 => n14998, A4 => 
                           n14997, ZN => n15018);
   U11865 : AND4_X1 port map( A1 => n14850, A2 => n14849, A3 => n14848, A4 => 
                           n14847, ZN => n14867);
   U11866 : AND4_X1 port map( A1 => n14678, A2 => n14677, A3 => n14676, A4 => 
                           n14675, ZN => n14695);
   U11867 : AND4_X1 port map( A1 => n14531, A2 => n14530, A3 => n14529, A4 => 
                           n14528, ZN => n14548);
   U11868 : AND4_X1 port map( A1 => n14380, A2 => n14379, A3 => n14378, A4 => 
                           n14377, ZN => n14397);
   U11869 : AND4_X1 port map( A1 => n14231, A2 => n14230, A3 => n14229, A4 => 
                           n14228, ZN => n14248);
   U11870 : AND4_X1 port map( A1 => n14083, A2 => n14082, A3 => n14081, A4 => 
                           n14080, ZN => n14100);
   U11871 : AND4_X1 port map( A1 => n13936, A2 => n13935, A3 => n13934, A4 => 
                           n13933, ZN => n13953);
   U11872 : AND4_X1 port map( A1 => n13789, A2 => n13788, A3 => n13787, A4 => 
                           n13786, ZN => n13806);
   U11873 : CLKBUF_X1 port map( A => n16797, Z => n16866);
   U11874 : CLKBUF_X1 port map( A => n16782, Z => n16851);
   U11875 : CLKBUF_X1 port map( A => n16767, Z => n16837);
   U11876 : CLKBUF_X1 port map( A => n16752, Z => n16822);
   U11877 : NAND2_X1 port map( A1 => n16678, A2 => n13731, ZN => n14910);
   U11878 : NAND3_X1 port map( A1 => ENABLE, A2 => RD1, A3 => n13731, ZN => 
                           n15166);
   U11879 : OR3_X2 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), A3 => n15166, 
                           ZN => n15115);
   U11880 : INV_X1 port map( A => ADD_RD1(2), ZN => n13733);
   U11881 : NAND3_X1 port map( A1 => n13733, A2 => n13734, A3 => ADD_RD1(1), ZN
                           => n13770);
   U11882 : NAND3_X1 port map( A1 => n13733, A2 => ADD_RD1(1), A3 => ADD_RD1(0)
                           , ZN => n13773);
   U11883 : CLKBUF_X2 port map( A => n15090, Z => n15121);
   U11884 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_63_port, B1 => 
                           n15121, B2 => REGISTERS_3_63_port, ZN => n13739);
   U11885 : INV_X1 port map( A => ADD_RD1(1), ZN => n13735);
   U11886 : NAND3_X1 port map( A1 => n13735, A2 => n13733, A3 => ADD_RD1(0), ZN
                           => n13768);
   U11887 : INV_X2 port map( A => n13768, ZN => n15065);
   U11888 : NAND2_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(0), ZN => n13732
                           );
   U11889 : INV_X2 port map( A => n13785, ZN => n15088);
   U11890 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_63_port, B1 => 
                           n15088, B2 => REGISTERS_5_63_port, ZN => n13738);
   U11891 : INV_X2 port map( A => n14461, ZN => n15091);
   U11892 : NAND3_X1 port map( A1 => n13735, A2 => n13733, A3 => n13734, ZN => 
                           n13756);
   U11893 : INV_X2 port map( A => n13756, ZN => n15089);
   U11894 : AOI22_X1 port map( A1 => n15091, A2 => REGISTERS_7_63_port, B1 => 
                           n15089, B2 => REGISTERS_0_63_port, ZN => n13737);
   U11895 : NAND3_X1 port map( A1 => n13734, A2 => ADD_RD1(2), A3 => ADD_RD1(1)
                           , ZN => n13771);
   U11896 : INV_X2 port map( A => n13771, ZN => n15043);
   U11897 : NAND3_X1 port map( A1 => n13735, A2 => n13734, A3 => ADD_RD1(2), ZN
                           => n13753);
   U11898 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_63_port, B1 => 
                           n15117, B2 => REGISTERS_4_63_port, ZN => n13736);
   U11899 : AND4_X1 port map( A1 => n13739, A2 => n13738, A3 => n13737, A4 => 
                           n13736, ZN => n13784);
   U11900 : CLKBUF_X2 port map( A => n15166, Z => n14354);
   U11901 : INV_X1 port map( A => ADD_RD1(4), ZN => n13742);
   U11902 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => n13742, ZN => n13766);
   U11903 : NOR2_X1 port map( A1 => n13766, A2 => n13773, ZN => n13740);
   U11904 : NOR2_X1 port map( A1 => n13766, A2 => n13753, ZN => n13741);
   U11905 : AOI22_X1 port map( A1 => REGISTERS_11_63_port, A2 => n15138, B1 => 
                           REGISTERS_12_63_port, B2 => n15140, ZN => n13752);
   U11906 : NOR2_X1 port map( A1 => n13772, A2 => n14461, ZN => n13743);
   U11907 : NOR2_X1 port map( A1 => n13772, A2 => n13753, ZN => n13744);
   U11908 : AOI22_X1 port map( A1 => REGISTERS_23_63_port, A2 => n15156, B1 => 
                           REGISTERS_20_63_port, B2 => n15153, ZN => n13751);
   U11909 : NOR2_X1 port map( A1 => n13766, A2 => n14461, ZN => n13745);
   U11910 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n13774
                           );
   U11911 : NOR2_X1 port map( A1 => n13774, A2 => n13756, ZN => n13746);
   U11912 : AOI22_X1 port map( A1 => REGISTERS_15_63_port, A2 => n15132, B1 => 
                           REGISTERS_24_63_port, B2 => n15127, ZN => n13750);
   U11913 : NOR2_X1 port map( A1 => n13772, A2 => n13756, ZN => n13747);
   U11914 : NOR2_X1 port map( A1 => n13774, A2 => n14461, ZN => n13748);
   U11915 : AOI22_X1 port map( A1 => REGISTERS_16_63_port, A2 => n15130, B1 => 
                           REGISTERS_31_63_port, B2 => n15152, ZN => n13749);
   U11916 : NAND4_X1 port map( A1 => n13752, A2 => n13751, A3 => n13750, A4 => 
                           n13749, ZN => n13782);
   U11917 : NOR2_X1 port map( A1 => n13774, A2 => n13753, ZN => n14837);
   U11918 : CLKBUF_X2 port map( A => n14837, Z => n15151);
   U11919 : NOR2_X1 port map( A1 => n13766, A2 => n13771, ZN => n13754);
   U11920 : AOI22_X1 port map( A1 => REGISTERS_28_63_port, A2 => n15151, B1 => 
                           REGISTERS_14_63_port, B2 => n15142, ZN => n13765);
   U11921 : NOR2_X1 port map( A1 => n13770, A2 => n13766, ZN => n13755);
   U11922 : NOR2_X1 port map( A1 => n13766, A2 => n13756, ZN => n13757);
   U11923 : AOI22_X1 port map( A1 => REGISTERS_10_63_port, A2 => n15150, B1 => 
                           REGISTERS_8_63_port, B2 => n15145, ZN => n13764);
   U11924 : NOR2_X1 port map( A1 => n13768, A2 => n13766, ZN => n13758);
   U11925 : NOR2_X1 port map( A1 => n13774, A2 => n13785, ZN => n13759);
   U11926 : AOI22_X1 port map( A1 => REGISTERS_9_63_port, A2 => n15144, B1 => 
                           REGISTERS_29_63_port, B2 => n15126, ZN => n13763);
   U11927 : NOR2_X1 port map( A1 => n13772, A2 => n13771, ZN => n13760);
   U11928 : NOR2_X1 port map( A1 => n13772, A2 => n13785, ZN => n13761);
   U11929 : AOI22_X1 port map( A1 => REGISTERS_22_63_port, A2 => n15128, B1 => 
                           REGISTERS_21_63_port, B2 => n15154, ZN => n13762);
   U11930 : NAND4_X1 port map( A1 => n13765, A2 => n13764, A3 => n13763, A4 => 
                           n13762, ZN => n13781);
   U11931 : NOR2_X1 port map( A1 => n13785, A2 => n13766, ZN => n13767);
   U11932 : NOR2_X1 port map( A1 => n13774, A2 => n13768, ZN => n14189);
   U11933 : AOI22_X1 port map( A1 => REGISTERS_13_63_port, A2 => n15157, B1 => 
                           REGISTERS_25_63_port, B2 => n14944, ZN => n13779);
   U11934 : NOR2_X1 port map( A1 => n13774, A2 => n13770, ZN => n15033);
   U11935 : NOR2_X1 port map( A1 => n13768, A2 => n13772, ZN => n13769);
   U11936 : AOI22_X1 port map( A1 => REGISTERS_26_63_port, A2 => n15033, B1 => 
                           REGISTERS_17_63_port, B2 => n15129, ZN => n13778);
   U11937 : NOR2_X1 port map( A1 => n13770, A2 => n13772, ZN => n14257);
   U11938 : CLKBUF_X2 port map( A => n14257, Z => n15101);
   U11939 : NOR2_X1 port map( A1 => n13774, A2 => n13771, ZN => n15032);
   U11940 : CLKBUF_X2 port map( A => n15032, Z => n15133);
   U11941 : AOI22_X1 port map( A1 => REGISTERS_18_63_port, A2 => n15101, B1 => 
                           REGISTERS_30_63_port, B2 => n15133, ZN => n13777);
   U11942 : NOR2_X1 port map( A1 => n13772, A2 => n13773, ZN => n14979);
   U11943 : NOR2_X1 port map( A1 => n13774, A2 => n13773, ZN => n13775);
   U11944 : AOI22_X1 port map( A1 => REGISTERS_19_63_port, A2 => n15139, B1 => 
                           REGISTERS_27_63_port, B2 => n15143, ZN => n13776);
   U11945 : NAND4_X1 port map( A1 => n13779, A2 => n13778, A3 => n13777, A4 => 
                           n13776, ZN => n13780);
   U11946 : NOR3_X1 port map( A1 => n13782, A2 => n13781, A3 => n13780, ZN => 
                           n13783);
   U11947 : OAI222_X1 port map( A1 => n16049, A2 => n8505, B1 => n15115, B2 => 
                           n13784, C1 => n14354, C2 => n13783, ZN => n8506);
   U11948 : CLKBUF_X2 port map( A => n15115, Z => n14505);
   U11949 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_62_port, B1 => 
                           n15091, B2 => REGISTERS_7_62_port, ZN => n13789);
   U11950 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_62_port, B1 => 
                           n15121, B2 => REGISTERS_3_62_port, ZN => n13788);
   U11951 : CLKBUF_X2 port map( A => n15117, Z => n14483);
   U11952 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_62_port, B1 => 
                           n14483, B2 => REGISTERS_4_62_port, ZN => n13787);
   U11953 : AOI22_X1 port map( A1 => n14781, A2 => REGISTERS_6_62_port, B1 => 
                           n15116, B2 => REGISTERS_0_62_port, ZN => n13786);
   U11954 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_62_port, B1 => 
                           n15150, B2 => REGISTERS_10_62_port, ZN => n13793);
   U11955 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_62_port, B1 => 
                           n15142, B2 => REGISTERS_14_62_port, ZN => n13792);
   U11956 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_62_port, B1 => 
                           n15154, B2 => REGISTERS_21_62_port, ZN => n13791);
   U11957 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_62_port, B1 => 
                           n15128, B2 => REGISTERS_22_62_port, ZN => n13790);
   U11958 : NAND4_X1 port map( A1 => n13793, A2 => n13792, A3 => n13791, A4 => 
                           n13790, ZN => n13804);
   U11959 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_62_port, B1 => 
                           n15145, B2 => REGISTERS_8_62_port, ZN => n13797);
   U11960 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_62_port, B1 => 
                           n15140, B2 => REGISTERS_12_62_port, ZN => n13796);
   U11961 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_62_port, B1 => 
                           n14837, B2 => REGISTERS_28_62_port, ZN => n13795);
   U11962 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_62_port, B1 => 
                           n15144, B2 => REGISTERS_9_62_port, ZN => n13794);
   U11963 : NAND4_X1 port map( A1 => n13797, A2 => n13796, A3 => n13795, A4 => 
                           n13794, ZN => n13803);
   U11964 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_62_port, B1 => 
                           n15130, B2 => REGISTERS_16_62_port, ZN => n13801);
   U11965 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_62_port, B1 => 
                           n15127, B2 => REGISTERS_24_62_port, ZN => n13800);
   U11966 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_62_port, B1 => 
                           n15138, B2 => REGISTERS_11_62_port, ZN => n13799);
   U11967 : CLKBUF_X2 port map( A => n15033, Z => n15131);
   U11968 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_62_port, B1 => 
                           n15126, B2 => REGISTERS_29_62_port, ZN => n13798);
   U11969 : NAND4_X1 port map( A1 => n13801, A2 => n13800, A3 => n13799, A4 => 
                           n13798, ZN => n13802);
   U11970 : NOR3_X1 port map( A1 => n13804, A2 => n13803, A3 => n13802, ZN => 
                           n13805);
   U11971 : OAI222_X1 port map( A1 => n16049, A2 => n8504, B1 => n14505, B2 => 
                           n13806, C1 => n15166, C2 => n13805, ZN => n8507);
   U11972 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_61_port, B1 => 
                           n15089, B2 => REGISTERS_0_61_port, ZN => n13810);
   U11973 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_61_port, B1 => 
                           n15091, B2 => REGISTERS_7_61_port, ZN => n13809);
   U11974 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_61_port, B1 => 
                           n15121, B2 => REGISTERS_3_61_port, ZN => n13808);
   U11975 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_61_port, B1 => 
                           n15117, B2 => REGISTERS_4_61_port, ZN => n13807);
   U11976 : AND4_X1 port map( A1 => n13810, A2 => n13809, A3 => n13808, A4 => 
                           n13807, ZN => n13827);
   U11977 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_61_port, B1 => 
                           n15142, B2 => REGISTERS_14_61_port, ZN => n13814);
   U11978 : AOI22_X1 port map( A1 => n15144, A2 => REGISTERS_9_61_port, B1 => 
                           n15126, B2 => REGISTERS_29_61_port, ZN => n13813);
   U11979 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_61_port, B1 => 
                           n15143, B2 => REGISTERS_27_61_port, ZN => n13812);
   U11980 : CLKBUF_X2 port map( A => n14189, Z => n14944);
   U11981 : AOI22_X1 port map( A1 => n15033, A2 => REGISTERS_26_61_port, B1 => 
                           n14944, B2 => REGISTERS_25_61_port, ZN => n13811);
   U11982 : NAND4_X1 port map( A1 => n13814, A2 => n13813, A3 => n13812, A4 => 
                           n13811, ZN => n13825);
   U11983 : CLKBUF_X2 port map( A => n14257, Z => n15155);
   U11984 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_61_port, B1 => 
                           n15153, B2 => REGISTERS_20_61_port, ZN => n13818);
   U11985 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_61_port, B1 => 
                           n15140, B2 => REGISTERS_12_61_port, ZN => n13817);
   U11986 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_61_port, B1 => 
                           n15150, B2 => REGISTERS_10_61_port, ZN => n13816);
   U11987 : AOI22_X1 port map( A1 => n15151, A2 => REGISTERS_28_61_port, B1 => 
                           n15128, B2 => REGISTERS_22_61_port, ZN => n13815);
   U11988 : NAND4_X1 port map( A1 => n13818, A2 => n13817, A3 => n13816, A4 => 
                           n13815, ZN => n13824);
   U11989 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_61_port, B1 => 
                           n15132, B2 => REGISTERS_15_61_port, ZN => n13822);
   U11990 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_61_port, B1 => 
                           n15145, B2 => REGISTERS_8_61_port, ZN => n13821);
   U11991 : CLKBUF_X2 port map( A => n14979, Z => n14832);
   U11992 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_61_port, B1 => 
                           n15130, B2 => REGISTERS_16_61_port, ZN => n13820);
   U11993 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_61_port, B1 => 
                           n15154, B2 => REGISTERS_21_61_port, ZN => n13819);
   U11994 : NAND4_X1 port map( A1 => n13822, A2 => n13821, A3 => n13820, A4 => 
                           n13819, ZN => n13823);
   U11995 : NOR3_X1 port map( A1 => n13825, A2 => n13824, A3 => n13823, ZN => 
                           n13826);
   U11996 : OAI222_X1 port map( A1 => n16049, A2 => n8503, B1 => n15115, B2 => 
                           n13827, C1 => n14354, C2 => n13826, ZN => n8508);
   U11997 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_60_port, B1 => 
                           n14483, B2 => REGISTERS_4_60_port, ZN => n13831);
   U11998 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_60_port, B1 => 
                           n15091, B2 => REGISTERS_7_60_port, ZN => n13830);
   U11999 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_60_port, B1 => 
                           n15121, B2 => REGISTERS_3_60_port, ZN => n13829);
   U12000 : AOI22_X1 port map( A1 => n14781, A2 => REGISTERS_6_60_port, B1 => 
                           n15116, B2 => REGISTERS_0_60_port, ZN => n13828);
   U12001 : AND4_X1 port map( A1 => n13831, A2 => n13830, A3 => n13829, A4 => 
                           n13828, ZN => n13848);
   U12002 : CLKBUF_X2 port map( A => n15032, Z => n15074);
   U12003 : AOI22_X1 port map( A1 => n15033, A2 => REGISTERS_26_60_port, B1 => 
                           n15074, B2 => REGISTERS_30_60_port, ZN => n13835);
   U12004 : AOI22_X1 port map( A1 => n15145, A2 => REGISTERS_8_60_port, B1 => 
                           n15154, B2 => REGISTERS_21_60_port, ZN => n13834);
   U12005 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_60_port, B1 => 
                           n15140, B2 => REGISTERS_12_60_port, ZN => n13833);
   U12006 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_60_port, B1 => 
                           n15096, B2 => REGISTERS_28_60_port, ZN => n13832);
   U12007 : NAND4_X1 port map( A1 => n13835, A2 => n13834, A3 => n13833, A4 => 
                           n13832, ZN => n13846);
   U12008 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_60_port, B1 => 
                           n15152, B2 => REGISTERS_31_60_port, ZN => n13839);
   U12009 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_60_port, B1 => 
                           n15138, B2 => REGISTERS_11_60_port, ZN => n13838);
   U12010 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_60_port, B1 => 
                           n15130, B2 => REGISTERS_16_60_port, ZN => n13837);
   U12011 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_60_port, B1 => 
                           n15150, B2 => REGISTERS_10_60_port, ZN => n13836);
   U12012 : NAND4_X1 port map( A1 => n13839, A2 => n13838, A3 => n13837, A4 => 
                           n13836, ZN => n13845);
   U12013 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_60_port, B1 => 
                           n15126, B2 => REGISTERS_29_60_port, ZN => n13843);
   U12014 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_60_port, B1 => 
                           n14979, B2 => REGISTERS_19_60_port, ZN => n13842);
   U12015 : AOI22_X1 port map( A1 => n15144, A2 => REGISTERS_9_60_port, B1 => 
                           n15128, B2 => REGISTERS_22_60_port, ZN => n13841);
   U12016 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_60_port, B1 => 
                           n15142, B2 => REGISTERS_14_60_port, ZN => n13840);
   U12017 : NAND4_X1 port map( A1 => n13843, A2 => n13842, A3 => n13841, A4 => 
                           n13840, ZN => n13844);
   U12018 : NOR3_X1 port map( A1 => n13846, A2 => n13845, A3 => n13844, ZN => 
                           n13847);
   U12019 : OAI222_X1 port map( A1 => n16049, A2 => n8502, B1 => n14505, B2 => 
                           n13848, C1 => n15166, C2 => n13847, ZN => n8509);
   U12020 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_59_port, B1 => 
                           n15117, B2 => REGISTERS_4_59_port, ZN => n13852);
   U12021 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_59_port, B1 => 
                           n15089, B2 => REGISTERS_0_59_port, ZN => n13851);
   U12022 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_59_port, B1 => 
                           n14781, B2 => REGISTERS_6_59_port, ZN => n13850);
   U12023 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_59_port, B1 => 
                           n15091, B2 => REGISTERS_7_59_port, ZN => n13849);
   U12024 : AND4_X1 port map( A1 => n13852, A2 => n13851, A3 => n13850, A4 => 
                           n13849, ZN => n13869);
   U12025 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_59_port, B1 => 
                           n15144, B2 => REGISTERS_9_59_port, ZN => n13856);
   U12026 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_59_port, B1 => 
                           n15145, B2 => REGISTERS_8_59_port, ZN => n13855);
   U12027 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_59_port, B1 => 
                           n15126, B2 => REGISTERS_29_59_port, ZN => n13854);
   U12028 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_59_port, B1 => 
                           n14944, B2 => REGISTERS_25_59_port, ZN => n13853);
   U12029 : NAND4_X1 port map( A1 => n13856, A2 => n13855, A3 => n13854, A4 => 
                           n13853, ZN => n13867);
   U12030 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_59_port, B1 => 
                           n15128, B2 => REGISTERS_22_59_port, ZN => n13860);
   U12031 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_59_port, B1 => 
                           n15142, B2 => REGISTERS_14_59_port, ZN => n13859);
   U12032 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_59_port, B1 => 
                           n15150, B2 => REGISTERS_10_59_port, ZN => n13858);
   U12033 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_59_port, B1 => 
                           n15101, B2 => REGISTERS_18_59_port, ZN => n13857);
   U12034 : NAND4_X1 port map( A1 => n13860, A2 => n13859, A3 => n13858, A4 => 
                           n13857, ZN => n13866);
   U12035 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_59_port, B1 => 
                           n15154, B2 => REGISTERS_21_59_port, ZN => n13864);
   U12036 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_59_port, B1 => 
                           n15140, B2 => REGISTERS_12_59_port, ZN => n13863);
   U12037 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_59_port, B1 => 
                           n15130, B2 => REGISTERS_16_59_port, ZN => n13862);
   U12038 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_59_port, B1 => 
                           n15151, B2 => REGISTERS_28_59_port, ZN => n13861);
   U12039 : NAND4_X1 port map( A1 => n13864, A2 => n13863, A3 => n13862, A4 => 
                           n13861, ZN => n13865);
   U12040 : NOR3_X1 port map( A1 => n13867, A2 => n13866, A3 => n13865, ZN => 
                           n13868);
   U12041 : OAI222_X1 port map( A1 => n16049, A2 => n8501, B1 => n14505, B2 => 
                           n13869, C1 => n14354, C2 => n13868, ZN => n8510);
   U12042 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_58_port, B1 => 
                           n14781, B2 => REGISTERS_6_58_port, ZN => n13873);
   U12043 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_58_port, B1 => 
                           n15121, B2 => REGISTERS_3_58_port, ZN => n13872);
   U12044 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_58_port, B1 => 
                           n15116, B2 => REGISTERS_0_58_port, ZN => n13871);
   U12045 : AOI22_X1 port map( A1 => n14483, A2 => REGISTERS_4_58_port, B1 => 
                           n15091, B2 => REGISTERS_7_58_port, ZN => n13870);
   U12046 : AND4_X1 port map( A1 => n13873, A2 => n13872, A3 => n13871, A4 => 
                           n13870, ZN => n13890);
   U12047 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_58_port, B1 => 
                           n15145, B2 => REGISTERS_8_58_port, ZN => n13877);
   U12048 : AOI22_X1 port map( A1 => n15126, A2 => REGISTERS_29_58_port, B1 => 
                           n15128, B2 => REGISTERS_22_58_port, ZN => n13876);
   U12049 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_58_port, B1 => 
                           n15127, B2 => REGISTERS_24_58_port, ZN => n13875);
   U12050 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_58_port, B1 => 
                           n15142, B2 => REGISTERS_14_58_port, ZN => n13874);
   U12051 : NAND4_X1 port map( A1 => n13877, A2 => n13876, A3 => n13875, A4 => 
                           n13874, ZN => n13888);
   U12052 : AOI22_X1 port map( A1 => n14979, A2 => REGISTERS_19_58_port, B1 => 
                           n15150, B2 => REGISTERS_10_58_port, ZN => n13881);
   U12053 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_58_port, B1 => 
                           n15132, B2 => REGISTERS_15_58_port, ZN => n13880);
   U12054 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_58_port, B1 => 
                           n15144, B2 => REGISTERS_9_58_port, ZN => n13879);
   U12055 : AOI22_X1 port map( A1 => n15033, A2 => REGISTERS_26_58_port, B1 => 
                           n15138, B2 => REGISTERS_11_58_port, ZN => n13878);
   U12056 : NAND4_X1 port map( A1 => n13881, A2 => n13880, A3 => n13879, A4 => 
                           n13878, ZN => n13887);
   U12057 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_58_port, B1 => 
                           n14837, B2 => REGISTERS_28_58_port, ZN => n13885);
   U12058 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_58_port, B1 => 
                           n15156, B2 => REGISTERS_23_58_port, ZN => n13884);
   U12059 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_58_port, B1 => 
                           n15153, B2 => REGISTERS_20_58_port, ZN => n13883);
   U12060 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_58_port, B1 => 
                           n15154, B2 => REGISTERS_21_58_port, ZN => n13882);
   U12061 : NAND4_X1 port map( A1 => n13885, A2 => n13884, A3 => n13883, A4 => 
                           n13882, ZN => n13886);
   U12062 : NOR3_X1 port map( A1 => n13888, A2 => n13887, A3 => n13886, ZN => 
                           n13889);
   U12063 : OAI222_X1 port map( A1 => n16049, A2 => n8500, B1 => n14505, B2 => 
                           n13890, C1 => n14354, C2 => n13889, ZN => n8511);
   U12064 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_57_port, B1 => 
                           n15091, B2 => REGISTERS_7_57_port, ZN => n13894);
   U12065 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_57_port, B1 => 
                           n14483, B2 => REGISTERS_4_57_port, ZN => n13893);
   U12066 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_57_port, B1 => 
                           n15043, B2 => REGISTERS_6_57_port, ZN => n13892);
   U12067 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_57_port, B1 => 
                           n15089, B2 => REGISTERS_0_57_port, ZN => n13891);
   U12068 : AND4_X1 port map( A1 => n13894, A2 => n13893, A3 => n13892, A4 => 
                           n13891, ZN => n13911);
   U12069 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_57_port, B1 => 
                           n15132, B2 => REGISTERS_15_57_port, ZN => n13898);
   U12070 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_57_port, B1 => 
                           n15145, B2 => REGISTERS_8_57_port, ZN => n13897);
   U12071 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_57_port, B1 => 
                           n15150, B2 => REGISTERS_10_57_port, ZN => n13896);
   U12072 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_57_port, B1 => 
                           n15128, B2 => REGISTERS_22_57_port, ZN => n13895);
   U12073 : NAND4_X1 port map( A1 => n13898, A2 => n13897, A3 => n13896, A4 => 
                           n13895, ZN => n13909);
   U12074 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_57_port, B1 => 
                           n15126, B2 => REGISTERS_29_57_port, ZN => n13902);
   U12075 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_57_port, B1 => 
                           n15127, B2 => REGISTERS_24_57_port, ZN => n13901);
   U12076 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_57_port, B1 => 
                           n15143, B2 => REGISTERS_27_57_port, ZN => n13900);
   U12077 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_57_port, B1 => 
                           n15142, B2 => REGISTERS_14_57_port, ZN => n13899);
   U12078 : NAND4_X1 port map( A1 => n13902, A2 => n13901, A3 => n13900, A4 => 
                           n13899, ZN => n13908);
   U12079 : AOI22_X1 port map( A1 => n14257, A2 => REGISTERS_18_57_port, B1 => 
                           n15096, B2 => REGISTERS_28_57_port, ZN => n13906);
   U12080 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_57_port, B1 => 
                           n15144, B2 => REGISTERS_9_57_port, ZN => n13905);
   U12081 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_57_port, B1 => 
                           n15152, B2 => REGISTERS_31_57_port, ZN => n13904);
   U12082 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_57_port, B1 => 
                           n15154, B2 => REGISTERS_21_57_port, ZN => n13903);
   U12083 : NAND4_X1 port map( A1 => n13906, A2 => n13905, A3 => n13904, A4 => 
                           n13903, ZN => n13907);
   U12084 : NOR3_X1 port map( A1 => n13909, A2 => n13908, A3 => n13907, ZN => 
                           n13910);
   U12085 : OAI222_X1 port map( A1 => n16049, A2 => n8499, B1 => n14505, B2 => 
                           n13911, C1 => n15166, C2 => n13910, ZN => n8512);
   U12086 : AOI22_X1 port map( A1 => n14781, A2 => REGISTERS_6_56_port, B1 => 
                           n15116, B2 => REGISTERS_0_56_port, ZN => n13915);
   U12087 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_56_port, B1 => 
                           n15091, B2 => REGISTERS_7_56_port, ZN => n13914);
   U12088 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_56_port, B1 => 
                           n15090, B2 => REGISTERS_3_56_port, ZN => n13913);
   U12089 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_56_port, B1 => 
                           n14483, B2 => REGISTERS_4_56_port, ZN => n13912);
   U12090 : AND4_X1 port map( A1 => n13915, A2 => n13914, A3 => n13913, A4 => 
                           n13912, ZN => n13932);
   U12091 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_56_port, B1 => 
                           n15128, B2 => REGISTERS_22_56_port, ZN => n13919);
   U12092 : AOI22_X1 port map( A1 => n14979, A2 => REGISTERS_19_56_port, B1 => 
                           n15154, B2 => REGISTERS_21_56_port, ZN => n13918);
   U12093 : AOI22_X1 port map( A1 => n15033, A2 => REGISTERS_26_56_port, B1 => 
                           n15150, B2 => REGISTERS_10_56_port, ZN => n13917);
   U12094 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_56_port, B1 => 
                           n15142, B2 => REGISTERS_14_56_port, ZN => n13916);
   U12095 : NAND4_X1 port map( A1 => n13919, A2 => n13918, A3 => n13917, A4 => 
                           n13916, ZN => n13930);
   U12096 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_56_port, B1 => 
                           n15144, B2 => REGISTERS_9_56_port, ZN => n13923);
   U12097 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_56_port, B1 => 
                           n15127, B2 => REGISTERS_24_56_port, ZN => n13922);
   U12098 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_56_port, B1 => 
                           n15101, B2 => REGISTERS_18_56_port, ZN => n13921);
   U12099 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_56_port, B1 => 
                           n15132, B2 => REGISTERS_15_56_port, ZN => n13920);
   U12100 : NAND4_X1 port map( A1 => n13923, A2 => n13922, A3 => n13921, A4 => 
                           n13920, ZN => n13929);
   U12101 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_56_port, B1 => 
                           n15151, B2 => REGISTERS_28_56_port, ZN => n13927);
   U12102 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_56_port, B1 => 
                           n15145, B2 => REGISTERS_8_56_port, ZN => n13926);
   U12103 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_56_port, B1 => 
                           n15126, B2 => REGISTERS_29_56_port, ZN => n13925);
   U12104 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_56_port, B1 => 
                           n15141, B2 => REGISTERS_25_56_port, ZN => n13924);
   U12105 : NAND4_X1 port map( A1 => n13927, A2 => n13926, A3 => n13925, A4 => 
                           n13924, ZN => n13928);
   U12106 : NOR3_X1 port map( A1 => n13930, A2 => n13929, A3 => n13928, ZN => 
                           n13931);
   U12107 : OAI222_X1 port map( A1 => n16049, A2 => n8498, B1 => n14505, B2 => 
                           n13932, C1 => n15166, C2 => n13931, ZN => n8513);
   U12108 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_55_port, B1 => 
                           n15091, B2 => REGISTERS_7_55_port, ZN => n13936);
   U12109 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_55_port, B1 => 
                           n15117, B2 => REGISTERS_4_55_port, ZN => n13935);
   U12110 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_55_port, B1 => 
                           n15089, B2 => REGISTERS_0_55_port, ZN => n13934);
   U12111 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_55_port, B1 => 
                           n15120, B2 => REGISTERS_1_55_port, ZN => n13933);
   U12112 : AOI22_X1 port map( A1 => n14979, A2 => REGISTERS_19_55_port, B1 => 
                           n15154, B2 => REGISTERS_21_55_port, ZN => n13940);
   U12113 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_55_port, B1 => 
                           n15153, B2 => REGISTERS_20_55_port, ZN => n13939);
   U12114 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_55_port, B1 => 
                           n15145, B2 => REGISTERS_8_55_port, ZN => n13938);
   U12115 : AOI22_X1 port map( A1 => n15151, A2 => REGISTERS_28_55_port, B1 => 
                           n15150, B2 => REGISTERS_10_55_port, ZN => n13937);
   U12116 : NAND4_X1 port map( A1 => n13940, A2 => n13939, A3 => n13938, A4 => 
                           n13937, ZN => n13951);
   U12117 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_55_port, B1 => 
                           n15126, B2 => REGISTERS_29_55_port, ZN => n13944);
   U12118 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_55_port, B1 => 
                           n15143, B2 => REGISTERS_27_55_port, ZN => n13943);
   U12119 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_55_port, B1 => 
                           n15142, B2 => REGISTERS_14_55_port, ZN => n13942);
   U12120 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_55_port, B1 => 
                           n15156, B2 => REGISTERS_23_55_port, ZN => n13941);
   U12121 : NAND4_X1 port map( A1 => n13944, A2 => n13943, A3 => n13942, A4 => 
                           n13941, ZN => n13950);
   U12122 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_55_port, B1 => 
                           n15130, B2 => REGISTERS_16_55_port, ZN => n13948);
   U12123 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_55_port, B1 => 
                           n15101, B2 => REGISTERS_18_55_port, ZN => n13947);
   U12124 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_55_port, B1 => 
                           n15144, B2 => REGISTERS_9_55_port, ZN => n13946);
   U12125 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_55_port, B1 => 
                           n15128, B2 => REGISTERS_22_55_port, ZN => n13945);
   U12126 : NAND4_X1 port map( A1 => n13948, A2 => n13947, A3 => n13946, A4 => 
                           n13945, ZN => n13949);
   U12127 : NOR3_X1 port map( A1 => n13951, A2 => n13950, A3 => n13949, ZN => 
                           n13952);
   U12128 : OAI222_X1 port map( A1 => n14910, A2 => n8497, B1 => n14505, B2 => 
                           n13953, C1 => n14354, C2 => n13952, ZN => n8514);
   U12129 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_54_port, B1 => 
                           n15121, B2 => REGISTERS_3_54_port, ZN => n13957);
   U12130 : AOI22_X1 port map( A1 => n14483, A2 => REGISTERS_4_54_port, B1 => 
                           n15091, B2 => REGISTERS_7_54_port, ZN => n13956);
   U12131 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_54_port, B1 => 
                           n14781, B2 => REGISTERS_6_54_port, ZN => n13955);
   U12132 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_54_port, B1 => 
                           n15116, B2 => REGISTERS_0_54_port, ZN => n13954);
   U12133 : AND4_X1 port map( A1 => n13957, A2 => n13956, A3 => n13955, A4 => 
                           n13954, ZN => n13974);
   U12134 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_54_port, B1 => 
                           n15145, B2 => REGISTERS_8_54_port, ZN => n13961);
   U12135 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_54_port, B1 => 
                           n15152, B2 => REGISTERS_31_54_port, ZN => n13960);
   U12136 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_54_port, B1 => 
                           n15142, B2 => REGISTERS_14_54_port, ZN => n13959);
   U12137 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_54_port, B1 => 
                           n15144, B2 => REGISTERS_9_54_port, ZN => n13958);
   U12138 : NAND4_X1 port map( A1 => n13961, A2 => n13960, A3 => n13959, A4 => 
                           n13958, ZN => n13972);
   U12139 : AOI22_X1 port map( A1 => n15033, A2 => REGISTERS_26_54_port, B1 => 
                           n15154, B2 => REGISTERS_21_54_port, ZN => n13965);
   U12140 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_54_port, B1 => 
                           n15138, B2 => REGISTERS_11_54_port, ZN => n13964);
   U12141 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_54_port, B1 => 
                           n15132, B2 => REGISTERS_15_54_port, ZN => n13963);
   U12142 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_54_port, B1 => 
                           n15153, B2 => REGISTERS_20_54_port, ZN => n13962);
   U12143 : NAND4_X1 port map( A1 => n13965, A2 => n13964, A3 => n13963, A4 => 
                           n13962, ZN => n13971);
   U12144 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_54_port, B1 => 
                           n14837, B2 => REGISTERS_28_54_port, ZN => n13969);
   U12145 : AOI22_X1 port map( A1 => n14257, A2 => REGISTERS_18_54_port, B1 => 
                           n15150, B2 => REGISTERS_10_54_port, ZN => n13968);
   U12146 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_54_port, B1 => 
                           n15128, B2 => REGISTERS_22_54_port, ZN => n13967);
   U12147 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_54_port, B1 => 
                           n15126, B2 => REGISTERS_29_54_port, ZN => n13966);
   U12148 : NAND4_X1 port map( A1 => n13969, A2 => n13968, A3 => n13967, A4 => 
                           n13966, ZN => n13970);
   U12149 : NOR3_X1 port map( A1 => n13972, A2 => n13971, A3 => n13970, ZN => 
                           n13973);
   U12150 : OAI222_X1 port map( A1 => n14910, A2 => n8496, B1 => n14505, B2 => 
                           n13974, C1 => n15166, C2 => n13973, ZN => n8515);
   U12151 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_53_port, B1 => 
                           n15117, B2 => REGISTERS_4_53_port, ZN => n13978);
   U12152 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_53_port, B1 => 
                           n15043, B2 => REGISTERS_6_53_port, ZN => n13977);
   U12153 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_53_port, B1 => 
                           n15089, B2 => REGISTERS_0_53_port, ZN => n13976);
   U12154 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_53_port, B1 => 
                           n15091, B2 => REGISTERS_7_53_port, ZN => n13975);
   U12155 : AND4_X1 port map( A1 => n13978, A2 => n13977, A3 => n13976, A4 => 
                           n13975, ZN => n13995);
   U12156 : AOI22_X1 port map( A1 => n15151, A2 => REGISTERS_28_53_port, B1 => 
                           n15144, B2 => REGISTERS_9_53_port, ZN => n13982);
   U12157 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_53_port, B1 => 
                           n15130, B2 => REGISTERS_16_53_port, ZN => n13981);
   U12158 : AOI22_X1 port map( A1 => n15128, A2 => REGISTERS_22_53_port, B1 => 
                           n15154, B2 => REGISTERS_21_53_port, ZN => n13980);
   U12159 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_53_port, B1 => 
                           n15150, B2 => REGISTERS_10_53_port, ZN => n13979);
   U12160 : NAND4_X1 port map( A1 => n13982, A2 => n13981, A3 => n13980, A4 => 
                           n13979, ZN => n13993);
   U12161 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_53_port, B1 => 
                           n15127, B2 => REGISTERS_24_53_port, ZN => n13986);
   U12162 : AOI22_X1 port map( A1 => n14979, A2 => REGISTERS_19_53_port, B1 => 
                           n15155, B2 => REGISTERS_18_53_port, ZN => n13985);
   U12163 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_53_port, B1 => 
                           n15156, B2 => REGISTERS_23_53_port, ZN => n13984);
   U12164 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_53_port, B1 => 
                           n15152, B2 => REGISTERS_31_53_port, ZN => n13983);
   U12165 : NAND4_X1 port map( A1 => n13986, A2 => n13985, A3 => n13984, A4 => 
                           n13983, ZN => n13992);
   U12166 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_53_port, B1 => 
                           n15145, B2 => REGISTERS_8_53_port, ZN => n13990);
   U12167 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_53_port, B1 => 
                           n15132, B2 => REGISTERS_15_53_port, ZN => n13989);
   U12168 : AOI22_X1 port map( A1 => n14189, A2 => REGISTERS_25_53_port, B1 => 
                           n15126, B2 => REGISTERS_29_53_port, ZN => n13988);
   U12169 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_53_port, B1 => 
                           n15142, B2 => REGISTERS_14_53_port, ZN => n13987);
   U12170 : NAND4_X1 port map( A1 => n13990, A2 => n13989, A3 => n13988, A4 => 
                           n13987, ZN => n13991);
   U12171 : NOR3_X1 port map( A1 => n13993, A2 => n13992, A3 => n13991, ZN => 
                           n13994);
   U12172 : OAI222_X1 port map( A1 => n14910, A2 => n8495, B1 => n14505, B2 => 
                           n13995, C1 => n14354, C2 => n13994, ZN => n8516);
   U12173 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_52_port, B1 => 
                           n15091, B2 => REGISTERS_7_52_port, ZN => n13999);
   U12174 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_52_port, B1 => 
                           n14781, B2 => REGISTERS_6_52_port, ZN => n13998);
   U12175 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_52_port, B1 => 
                           n15116, B2 => REGISTERS_0_52_port, ZN => n13997);
   U12176 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_52_port, B1 => 
                           n14483, B2 => REGISTERS_4_52_port, ZN => n13996);
   U12177 : AND4_X1 port map( A1 => n13999, A2 => n13998, A3 => n13997, A4 => 
                           n13996, ZN => n14016);
   U12178 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_52_port, B1 => 
                           n15154, B2 => REGISTERS_21_52_port, ZN => n14003);
   U12179 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_52_port, B1 => 
                           n15140, B2 => REGISTERS_12_52_port, ZN => n14002);
   U12180 : AOI22_X1 port map( A1 => n15033, A2 => REGISTERS_26_52_port, B1 => 
                           n15142, B2 => REGISTERS_14_52_port, ZN => n14001);
   U12181 : AOI22_X1 port map( A1 => n14189, A2 => REGISTERS_25_52_port, B1 => 
                           n15074, B2 => REGISTERS_30_52_port, ZN => n14000);
   U12182 : NAND4_X1 port map( A1 => n14003, A2 => n14002, A3 => n14001, A4 => 
                           n14000, ZN => n14014);
   U12183 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_52_port, B1 => 
                           n15151, B2 => REGISTERS_28_52_port, ZN => n14007);
   U12184 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_52_port, B1 => 
                           n15145, B2 => REGISTERS_8_52_port, ZN => n14006);
   U12185 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_52_port, B1 => 
                           n15153, B2 => REGISTERS_20_52_port, ZN => n14005);
   U12186 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_52_port, B1 => 
                           n15138, B2 => REGISTERS_11_52_port, ZN => n14004);
   U12187 : NAND4_X1 port map( A1 => n14007, A2 => n14006, A3 => n14005, A4 => 
                           n14004, ZN => n14013);
   U12188 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_52_port, B1 => 
                           n15127, B2 => REGISTERS_24_52_port, ZN => n14011);
   U12189 : AOI22_X1 port map( A1 => n15144, A2 => REGISTERS_9_52_port, B1 => 
                           n15128, B2 => REGISTERS_22_52_port, ZN => n14010);
   U12190 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_52_port, B1 => 
                           n15126, B2 => REGISTERS_29_52_port, ZN => n14009);
   U12191 : AOI22_X1 port map( A1 => n14257, A2 => REGISTERS_18_52_port, B1 => 
                           n15130, B2 => REGISTERS_16_52_port, ZN => n14008);
   U12192 : NAND4_X1 port map( A1 => n14011, A2 => n14010, A3 => n14009, A4 => 
                           n14008, ZN => n14012);
   U12193 : NOR3_X1 port map( A1 => n14014, A2 => n14013, A3 => n14012, ZN => 
                           n14015);
   U12194 : OAI222_X1 port map( A1 => n14910, A2 => n8494, B1 => n14505, B2 => 
                           n14016, C1 => n15166, C2 => n14015, ZN => n8517);
   U12195 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_51_port, B1 => 
                           n14781, B2 => REGISTERS_6_51_port, ZN => n14020);
   U12196 : AOI22_X1 port map( A1 => n15091, A2 => REGISTERS_7_51_port, B1 => 
                           n15089, B2 => REGISTERS_0_51_port, ZN => n14019);
   U12197 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_51_port, B1 => 
                           n15088, B2 => REGISTERS_5_51_port, ZN => n14018);
   U12198 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_51_port, B1 => 
                           n15117, B2 => REGISTERS_4_51_port, ZN => n14017);
   U12199 : AND4_X1 port map( A1 => n14020, A2 => n14019, A3 => n14018, A4 => 
                           n14017, ZN => n14037);
   U12200 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_51_port, B1 => 
                           n15145, B2 => REGISTERS_8_51_port, ZN => n14024);
   U12201 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_51_port, B1 => 
                           n15130, B2 => REGISTERS_16_51_port, ZN => n14023);
   U12202 : CLKBUF_X2 port map( A => n15131, Z => n15005);
   U12203 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_51_port, B1 => 
                           n15127, B2 => REGISTERS_24_51_port, ZN => n14022);
   U12204 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_51_port, B1 => 
                           n15150, B2 => REGISTERS_10_51_port, ZN => n14021);
   U12205 : NAND4_X1 port map( A1 => n14024, A2 => n14023, A3 => n14022, A4 => 
                           n14021, ZN => n14035);
   U12206 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_51_port, B1 => 
                           n15144, B2 => REGISTERS_9_51_port, ZN => n14028);
   U12207 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_51_port, B1 => 
                           n15154, B2 => REGISTERS_21_51_port, ZN => n14027);
   U12208 : AOI22_X1 port map( A1 => n15126, A2 => REGISTERS_29_51_port, B1 => 
                           n15128, B2 => REGISTERS_22_51_port, ZN => n14026);
   U12209 : AOI22_X1 port map( A1 => n14189, A2 => REGISTERS_25_51_port, B1 => 
                           n15143, B2 => REGISTERS_27_51_port, ZN => n14025);
   U12210 : NAND4_X1 port map( A1 => n14028, A2 => n14027, A3 => n14026, A4 => 
                           n14025, ZN => n14034);
   U12211 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_51_port, B1 => 
                           n15138, B2 => REGISTERS_11_51_port, ZN => n14032);
   U12212 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_51_port, B1 => 
                           n15156, B2 => REGISTERS_23_51_port, ZN => n14031);
   U12213 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_51_port, B1 => 
                           n15096, B2 => REGISTERS_28_51_port, ZN => n14030);
   U12214 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_51_port, B1 => 
                           n15142, B2 => REGISTERS_14_51_port, ZN => n14029);
   U12215 : NAND4_X1 port map( A1 => n14032, A2 => n14031, A3 => n14030, A4 => 
                           n14029, ZN => n14033);
   U12216 : NOR3_X1 port map( A1 => n14035, A2 => n14034, A3 => n14033, ZN => 
                           n14036);
   U12217 : OAI222_X1 port map( A1 => n14910, A2 => n8493, B1 => n15115, B2 => 
                           n14037, C1 => n14354, C2 => n14036, ZN => n8518);
   U12218 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_50_port, B1 => 
                           n15121, B2 => REGISTERS_3_50_port, ZN => n14041);
   U12219 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_50_port, B1 => 
                           n15091, B2 => REGISTERS_7_50_port, ZN => n14040);
   U12220 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_50_port, B1 => 
                           n14483, B2 => REGISTERS_4_50_port, ZN => n14039);
   U12221 : AOI22_X1 port map( A1 => n14781, A2 => REGISTERS_6_50_port, B1 => 
                           n15089, B2 => REGISTERS_0_50_port, ZN => n14038);
   U12222 : AND4_X1 port map( A1 => n14041, A2 => n14040, A3 => n14039, A4 => 
                           n14038, ZN => n14058);
   U12223 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_50_port, B1 => 
                           n15096, B2 => REGISTERS_28_50_port, ZN => n14045);
   U12224 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_50_port, B1 => 
                           n15127, B2 => REGISTERS_24_50_port, ZN => n14044);
   U12225 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_50_port, B1 => 
                           n15126, B2 => REGISTERS_29_50_port, ZN => n14043);
   U12226 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_50_port, B1 => 
                           n15145, B2 => REGISTERS_8_50_port, ZN => n14042);
   U12227 : NAND4_X1 port map( A1 => n14045, A2 => n14044, A3 => n14043, A4 => 
                           n14042, ZN => n14056);
   U12228 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_50_port, B1 => 
                           n15154, B2 => REGISTERS_21_50_port, ZN => n14049);
   U12229 : AOI22_X1 port map( A1 => n14189, A2 => REGISTERS_25_50_port, B1 => 
                           n15128, B2 => REGISTERS_22_50_port, ZN => n14048);
   U12230 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_50_port, B1 => 
                           n15142, B2 => REGISTERS_14_50_port, ZN => n14047);
   U12231 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_50_port, B1 => 
                           n15152, B2 => REGISTERS_31_50_port, ZN => n14046);
   U12232 : NAND4_X1 port map( A1 => n14049, A2 => n14048, A3 => n14047, A4 => 
                           n14046, ZN => n14055);
   U12233 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_50_port, B1 => 
                           n15130, B2 => REGISTERS_16_50_port, ZN => n14053);
   U12234 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_50_port, B1 => 
                           n15150, B2 => REGISTERS_10_50_port, ZN => n14052);
   U12235 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_50_port, B1 => 
                           n15144, B2 => REGISTERS_9_50_port, ZN => n14051);
   U12236 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_50_port, B1 => 
                           n15132, B2 => REGISTERS_15_50_port, ZN => n14050);
   U12237 : NAND4_X1 port map( A1 => n14053, A2 => n14052, A3 => n14051, A4 => 
                           n14050, ZN => n14054);
   U12238 : NOR3_X1 port map( A1 => n14056, A2 => n14055, A3 => n14054, ZN => 
                           n14057);
   U12239 : OAI222_X1 port map( A1 => n14910, A2 => n8492, B1 => n14505, B2 => 
                           n14058, C1 => n14354, C2 => n14057, ZN => n8519);
   U12240 : CLKBUF_X2 port map( A => n14910, Z => n16071);
   U12241 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_49_port, B1 => 
                           n15091, B2 => REGISTERS_7_49_port, ZN => n14062);
   U12242 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_49_port, B1 => 
                           n15089, B2 => REGISTERS_0_49_port, ZN => n14061);
   U12243 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_49_port, B1 => 
                           n15090, B2 => REGISTERS_3_49_port, ZN => n14060);
   U12244 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_49_port, B1 => 
                           n15117, B2 => REGISTERS_4_49_port, ZN => n14059);
   U12245 : AND4_X1 port map( A1 => n14062, A2 => n14061, A3 => n14060, A4 => 
                           n14059, ZN => n14079);
   U12246 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_49_port, B1 => 
                           n15138, B2 => REGISTERS_11_49_port, ZN => n14066);
   U12247 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_49_port, B1 => 
                           n15151, B2 => REGISTERS_28_49_port, ZN => n14065);
   U12248 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_49_port, B1 => 
                           n14979, B2 => REGISTERS_19_49_port, ZN => n14064);
   U12249 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_49_port, B1 => 
                           n15144, B2 => REGISTERS_9_49_port, ZN => n14063);
   U12250 : NAND4_X1 port map( A1 => n14066, A2 => n14065, A3 => n14064, A4 => 
                           n14063, ZN => n14077);
   U12251 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_49_port, B1 => 
                           n15154, B2 => REGISTERS_21_49_port, ZN => n14070);
   U12252 : AOI22_X1 port map( A1 => n15142, A2 => REGISTERS_14_49_port, B1 => 
                           n15150, B2 => REGISTERS_10_49_port, ZN => n14069);
   U12253 : AOI22_X1 port map( A1 => n14257, A2 => REGISTERS_18_49_port, B1 => 
                           n15140, B2 => REGISTERS_12_49_port, ZN => n14068);
   U12254 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_49_port, B1 => 
                           n15128, B2 => REGISTERS_22_49_port, ZN => n14067);
   U12255 : NAND4_X1 port map( A1 => n14070, A2 => n14069, A3 => n14068, A4 => 
                           n14067, ZN => n14076);
   U12256 : AOI22_X1 port map( A1 => n14189, A2 => REGISTERS_25_49_port, B1 => 
                           n15156, B2 => REGISTERS_23_49_port, ZN => n14074);
   U12257 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_49_port, B1 => 
                           n15152, B2 => REGISTERS_31_49_port, ZN => n14073);
   U12258 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_49_port, B1 => 
                           n15145, B2 => REGISTERS_8_49_port, ZN => n14072);
   U12259 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_49_port, B1 => 
                           n15126, B2 => REGISTERS_29_49_port, ZN => n14071);
   U12260 : NAND4_X1 port map( A1 => n14074, A2 => n14073, A3 => n14072, A4 => 
                           n14071, ZN => n14075);
   U12261 : NOR3_X1 port map( A1 => n14077, A2 => n14076, A3 => n14075, ZN => 
                           n14078);
   U12262 : OAI222_X1 port map( A1 => n16071, A2 => n8491, B1 => n14505, B2 => 
                           n14079, C1 => n15166, C2 => n14078, ZN => n8520);
   U12263 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_48_port, B1 => 
                           n15089, B2 => REGISTERS_0_48_port, ZN => n14083);
   U12264 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_48_port, B1 => 
                           n15121, B2 => REGISTERS_3_48_port, ZN => n14082);
   U12265 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_48_port, B1 => 
                           n14483, B2 => REGISTERS_4_48_port, ZN => n14081);
   U12266 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_48_port, B1 => 
                           n15091, B2 => REGISTERS_7_48_port, ZN => n14080);
   U12267 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_48_port, B1 => 
                           n15128, B2 => REGISTERS_22_48_port, ZN => n14087);
   U12268 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_48_port, B1 => 
                           n15150, B2 => REGISTERS_10_48_port, ZN => n14086);
   U12269 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_48_port, B1 => 
                           n15156, B2 => REGISTERS_23_48_port, ZN => n14085);
   U12270 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_48_port, B1 => 
                           n15126, B2 => REGISTERS_29_48_port, ZN => n14084);
   U12271 : NAND4_X1 port map( A1 => n14087, A2 => n14086, A3 => n14085, A4 => 
                           n14084, ZN => n14098);
   U12272 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_48_port, B1 => 
                           n15127, B2 => REGISTERS_24_48_port, ZN => n14091);
   U12273 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_48_port, B1 => 
                           n15144, B2 => REGISTERS_9_48_port, ZN => n14090);
   U12274 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_48_port, B1 => 
                           n15130, B2 => REGISTERS_16_48_port, ZN => n14089);
   U12275 : CLKBUF_X2 port map( A => n14979, Z => n15139);
   U12276 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_48_port, B1 => 
                           n15154, B2 => REGISTERS_21_48_port, ZN => n14088);
   U12277 : NAND4_X1 port map( A1 => n14091, A2 => n14090, A3 => n14089, A4 => 
                           n14088, ZN => n14097);
   U12278 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_48_port, B1 => 
                           n15101, B2 => REGISTERS_18_48_port, ZN => n14095);
   U12279 : AOI22_X1 port map( A1 => n15151, A2 => REGISTERS_28_48_port, B1 => 
                           n15142, B2 => REGISTERS_14_48_port, ZN => n14094);
   U12280 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_48_port, B1 => 
                           n15153, B2 => REGISTERS_20_48_port, ZN => n14093);
   U12281 : AOI22_X1 port map( A1 => n14189, A2 => REGISTERS_25_48_port, B1 => 
                           n15145, B2 => REGISTERS_8_48_port, ZN => n14092);
   U12282 : NAND4_X1 port map( A1 => n14095, A2 => n14094, A3 => n14093, A4 => 
                           n14092, ZN => n14096);
   U12283 : NOR3_X1 port map( A1 => n14098, A2 => n14097, A3 => n14096, ZN => 
                           n14099);
   U12284 : OAI222_X1 port map( A1 => n14910, A2 => n8490, B1 => n15115, B2 => 
                           n14100, C1 => n15166, C2 => n14099, ZN => n8521);
   U12285 : AOI22_X1 port map( A1 => n15117, A2 => REGISTERS_4_47_port, B1 => 
                           n15089, B2 => REGISTERS_0_47_port, ZN => n14104);
   U12286 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_47_port, B1 => 
                           n15121, B2 => REGISTERS_3_47_port, ZN => n14103);
   U12287 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_47_port, B1 => 
                           n15119, B2 => REGISTERS_7_47_port, ZN => n14102);
   U12288 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_47_port, B1 => 
                           n15043, B2 => REGISTERS_6_47_port, ZN => n14101);
   U12289 : AND4_X1 port map( A1 => n14104, A2 => n14103, A3 => n14102, A4 => 
                           n14101, ZN => n14121);
   U12290 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_47_port, B1 => 
                           n15154, B2 => REGISTERS_21_47_port, ZN => n14108);
   U12291 : AOI22_X1 port map( A1 => n14189, A2 => REGISTERS_25_47_port, B1 => 
                           n15142, B2 => REGISTERS_14_47_port, ZN => n14107);
   U12292 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_47_port, B1 => 
                           n15032, B2 => REGISTERS_30_47_port, ZN => n14106);
   U12293 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_47_port, B1 => 
                           n15144, B2 => REGISTERS_9_47_port, ZN => n14105);
   U12294 : NAND4_X1 port map( A1 => n14108, A2 => n14107, A3 => n14106, A4 => 
                           n14105, ZN => n14119);
   U12295 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_47_port, B1 => 
                           n15151, B2 => REGISTERS_28_47_port, ZN => n14112);
   U12296 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_47_port, B1 => 
                           n15126, B2 => REGISTERS_29_47_port, ZN => n14111);
   U12297 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_47_port, B1 => 
                           n15152, B2 => REGISTERS_31_47_port, ZN => n14110);
   U12298 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_47_port, B1 => 
                           n15140, B2 => REGISTERS_12_47_port, ZN => n14109);
   U12299 : NAND4_X1 port map( A1 => n14112, A2 => n14111, A3 => n14110, A4 => 
                           n14109, ZN => n14118);
   U12300 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_47_port, B1 => 
                           n15127, B2 => REGISTERS_24_47_port, ZN => n14116);
   U12301 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_47_port, B1 => 
                           n15155, B2 => REGISTERS_18_47_port, ZN => n14115);
   U12302 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_47_port, B1 => 
                           n15128, B2 => REGISTERS_22_47_port, ZN => n14114);
   U12303 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_47_port, B1 => 
                           n15145, B2 => REGISTERS_8_47_port, ZN => n14113);
   U12304 : NAND4_X1 port map( A1 => n14116, A2 => n14115, A3 => n14114, A4 => 
                           n14113, ZN => n14117);
   U12305 : NOR3_X1 port map( A1 => n14119, A2 => n14118, A3 => n14117, ZN => 
                           n14120);
   U12306 : OAI222_X1 port map( A1 => n16071, A2 => n8489, B1 => n15115, B2 => 
                           n14121, C1 => n14354, C2 => n14120, ZN => n8522);
   U12307 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_46_port, B1 => 
                           n15043, B2 => REGISTERS_6_46_port, ZN => n14125);
   U12308 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_46_port, B1 => 
                           n15121, B2 => REGISTERS_3_46_port, ZN => n14124);
   U12309 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_46_port, B1 => 
                           n14483, B2 => REGISTERS_4_46_port, ZN => n14123);
   U12310 : AOI22_X1 port map( A1 => n15091, A2 => REGISTERS_7_46_port, B1 => 
                           n15089, B2 => REGISTERS_0_46_port, ZN => n14122);
   U12311 : AND4_X1 port map( A1 => n14125, A2 => n14124, A3 => n14123, A4 => 
                           n14122, ZN => n14142);
   U12312 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_46_port, B1 => 
                           n15153, B2 => REGISTERS_20_46_port, ZN => n14129);
   U12313 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_46_port, B1 => 
                           n15140, B2 => REGISTERS_12_46_port, ZN => n14128);
   U12314 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_46_port, B1 => 
                           n15145, B2 => REGISTERS_8_46_port, ZN => n14127);
   U12315 : AOI22_X1 port map( A1 => n14257, A2 => REGISTERS_18_46_port, B1 => 
                           n15128, B2 => REGISTERS_22_46_port, ZN => n14126);
   U12316 : NAND4_X1 port map( A1 => n14129, A2 => n14128, A3 => n14127, A4 => 
                           n14126, ZN => n14140);
   U12317 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_46_port, B1 => 
                           n15152, B2 => REGISTERS_31_46_port, ZN => n14133);
   U12318 : AOI22_X1 port map( A1 => n14189, A2 => REGISTERS_25_46_port, B1 => 
                           n15126, B2 => REGISTERS_29_46_port, ZN => n14132);
   U12319 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_46_port, B1 => 
                           n15032, B2 => REGISTERS_30_46_port, ZN => n14131);
   U12320 : AOI22_X1 port map( A1 => n15151, A2 => REGISTERS_28_46_port, B1 => 
                           n15142, B2 => REGISTERS_14_46_port, ZN => n14130);
   U12321 : NAND4_X1 port map( A1 => n14133, A2 => n14132, A3 => n14131, A4 => 
                           n14130, ZN => n14139);
   U12322 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_46_port, B1 => 
                           n15154, B2 => REGISTERS_21_46_port, ZN => n14137);
   U12323 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_46_port, B1 => 
                           n15144, B2 => REGISTERS_9_46_port, ZN => n14136);
   U12324 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_46_port, B1 => 
                           n15143, B2 => REGISTERS_27_46_port, ZN => n14135);
   U12325 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_46_port, B1 => 
                           n15127, B2 => REGISTERS_24_46_port, ZN => n14134);
   U12326 : NAND4_X1 port map( A1 => n14137, A2 => n14136, A3 => n14135, A4 => 
                           n14134, ZN => n14138);
   U12327 : NOR3_X1 port map( A1 => n14140, A2 => n14139, A3 => n14138, ZN => 
                           n14141);
   U12328 : OAI222_X1 port map( A1 => n14910, A2 => n8488, B1 => n14505, B2 => 
                           n14142, C1 => n14354, C2 => n14141, ZN => n8523);
   U12329 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_45_port, B1 => 
                           n15121, B2 => REGISTERS_3_45_port, ZN => n14146);
   U12330 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_45_port, B1 => 
                           n15089, B2 => REGISTERS_0_45_port, ZN => n14145);
   U12331 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_45_port, B1 => 
                           n15091, B2 => REGISTERS_7_45_port, ZN => n14144);
   U12332 : AOI22_X1 port map( A1 => n14781, A2 => REGISTERS_6_45_port, B1 => 
                           n15117, B2 => REGISTERS_4_45_port, ZN => n14143);
   U12333 : AND4_X1 port map( A1 => n14146, A2 => n14145, A3 => n14144, A4 => 
                           n14143, ZN => n14163);
   U12334 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_45_port, B1 => 
                           n15142, B2 => REGISTERS_14_45_port, ZN => n14150);
   U12335 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_45_port, B1 => 
                           n15156, B2 => REGISTERS_23_45_port, ZN => n14149);
   U12336 : AOI22_X1 port map( A1 => n14189, A2 => REGISTERS_25_45_port, B1 => 
                           n15150, B2 => REGISTERS_10_45_port, ZN => n14148);
   U12337 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_45_port, B1 => 
                           n15154, B2 => REGISTERS_21_45_port, ZN => n14147);
   U12338 : NAND4_X1 port map( A1 => n14150, A2 => n14149, A3 => n14148, A4 => 
                           n14147, ZN => n14161);
   U12339 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_45_port, B1 => 
                           n15143, B2 => REGISTERS_27_45_port, ZN => n14154);
   U12340 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_45_port, B1 => 
                           n15132, B2 => REGISTERS_15_45_port, ZN => n14153);
   U12341 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_45_port, B1 => 
                           n15152, B2 => REGISTERS_31_45_port, ZN => n14152);
   U12342 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_45_port, B1 => 
                           n15153, B2 => REGISTERS_20_45_port, ZN => n14151);
   U12343 : NAND4_X1 port map( A1 => n14154, A2 => n14153, A3 => n14152, A4 => 
                           n14151, ZN => n14160);
   U12344 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_45_port, B1 => 
                           n15128, B2 => REGISTERS_22_45_port, ZN => n14158);
   U12345 : AOI22_X1 port map( A1 => n14257, A2 => REGISTERS_18_45_port, B1 => 
                           n15145, B2 => REGISTERS_8_45_port, ZN => n14157);
   U12346 : AOI22_X1 port map( A1 => n15151, A2 => REGISTERS_28_45_port, B1 => 
                           n15126, B2 => REGISTERS_29_45_port, ZN => n14156);
   U12347 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_45_port, B1 => 
                           n15144, B2 => REGISTERS_9_45_port, ZN => n14155);
   U12348 : NAND4_X1 port map( A1 => n14158, A2 => n14157, A3 => n14156, A4 => 
                           n14155, ZN => n14159);
   U12349 : NOR3_X1 port map( A1 => n14161, A2 => n14160, A3 => n14159, ZN => 
                           n14162);
   U12350 : OAI222_X1 port map( A1 => n16071, A2 => n8487, B1 => n14505, B2 => 
                           n14163, C1 => n14354, C2 => n14162, ZN => n8524);
   U12351 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_44_port, B1 => 
                           n15088, B2 => REGISTERS_5_44_port, ZN => n14167);
   U12352 : AOI22_X1 port map( A1 => n15091, A2 => REGISTERS_7_44_port, B1 => 
                           n15089, B2 => REGISTERS_0_44_port, ZN => n14166);
   U12353 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_44_port, B1 => 
                           n15117, B2 => REGISTERS_4_44_port, ZN => n14165);
   U12354 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_44_port, B1 => 
                           n14781, B2 => REGISTERS_6_44_port, ZN => n14164);
   U12355 : AND4_X1 port map( A1 => n14167, A2 => n14166, A3 => n14165, A4 => 
                           n14164, ZN => n14184);
   U12356 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_44_port, B1 => 
                           n15130, B2 => REGISTERS_16_44_port, ZN => n14171);
   U12357 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_44_port, B1 => 
                           n15154, B2 => REGISTERS_21_44_port, ZN => n14170);
   U12358 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_44_port, B1 => 
                           n15132, B2 => REGISTERS_15_44_port, ZN => n14169);
   U12359 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_44_port, B1 => 
                           n15128, B2 => REGISTERS_22_44_port, ZN => n14168);
   U12360 : NAND4_X1 port map( A1 => n14171, A2 => n14170, A3 => n14169, A4 => 
                           n14168, ZN => n14182);
   U12361 : AOI22_X1 port map( A1 => n15145, A2 => REGISTERS_8_44_port, B1 => 
                           n15126, B2 => REGISTERS_29_44_port, ZN => n14175);
   U12362 : AOI22_X1 port map( A1 => n14257, A2 => REGISTERS_18_44_port, B1 => 
                           n15127, B2 => REGISTERS_24_44_port, ZN => n14174);
   U12363 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_44_port, B1 => 
                           n15142, B2 => REGISTERS_14_44_port, ZN => n14173);
   U12364 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_44_port, B1 => 
                           n15138, B2 => REGISTERS_11_44_port, ZN => n14172);
   U12365 : NAND4_X1 port map( A1 => n14175, A2 => n14174, A3 => n14173, A4 => 
                           n14172, ZN => n14181);
   U12366 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_44_port, B1 => 
                           n15144, B2 => REGISTERS_9_44_port, ZN => n14179);
   U12367 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_44_port, B1 => 
                           n15139, B2 => REGISTERS_19_44_port, ZN => n14178);
   U12368 : AOI22_X1 port map( A1 => n14189, A2 => REGISTERS_25_44_port, B1 => 
                           n15152, B2 => REGISTERS_31_44_port, ZN => n14177);
   U12369 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_44_port, B1 => 
                           n15096, B2 => REGISTERS_28_44_port, ZN => n14176);
   U12370 : NAND4_X1 port map( A1 => n14179, A2 => n14178, A3 => n14177, A4 => 
                           n14176, ZN => n14180);
   U12371 : NOR3_X1 port map( A1 => n14182, A2 => n14181, A3 => n14180, ZN => 
                           n14183);
   U12372 : OAI222_X1 port map( A1 => n14910, A2 => n8486, B1 => n15115, B2 => 
                           n14184, C1 => n14354, C2 => n14183, ZN => n8525);
   U12373 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_43_port, B1 => 
                           n15089, B2 => REGISTERS_0_43_port, ZN => n14188);
   U12374 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_43_port, B1 => 
                           n15119, B2 => REGISTERS_7_43_port, ZN => n14187);
   U12375 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_43_port, B1 => 
                           n15088, B2 => REGISTERS_5_43_port, ZN => n14186);
   U12376 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_43_port, B1 => 
                           n14483, B2 => REGISTERS_4_43_port, ZN => n14185);
   U12377 : AND4_X1 port map( A1 => n14188, A2 => n14187, A3 => n14186, A4 => 
                           n14185, ZN => n14206);
   U12378 : AOI22_X1 port map( A1 => n15142, A2 => REGISTERS_14_43_port, B1 => 
                           n15145, B2 => REGISTERS_8_43_port, ZN => n14193);
   U12379 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_43_port, B1 => 
                           n15150, B2 => REGISTERS_10_43_port, ZN => n14192);
   U12380 : CLKBUF_X2 port map( A => n14189, Z => n15141);
   U12381 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_43_port, B1 => 
                           n15153, B2 => REGISTERS_20_43_port, ZN => n14191);
   U12382 : AOI22_X1 port map( A1 => n14257, A2 => REGISTERS_18_43_port, B1 => 
                           n15154, B2 => REGISTERS_21_43_port, ZN => n14190);
   U12383 : NAND4_X1 port map( A1 => n14193, A2 => n14192, A3 => n14191, A4 => 
                           n14190, ZN => n14204);
   U12384 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_43_port, B1 => 
                           n15143, B2 => REGISTERS_27_43_port, ZN => n14197);
   U12385 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_43_port, B1 => 
                           n15152, B2 => REGISTERS_31_43_port, ZN => n14196);
   U12386 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_43_port, B1 => 
                           n15128, B2 => REGISTERS_22_43_port, ZN => n14195);
   U12387 : AOI22_X1 port map( A1 => n15151, A2 => REGISTERS_28_43_port, B1 => 
                           n15126, B2 => REGISTERS_29_43_port, ZN => n14194);
   U12388 : NAND4_X1 port map( A1 => n14197, A2 => n14196, A3 => n14195, A4 => 
                           n14194, ZN => n14203);
   U12389 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_43_port, B1 => 
                           n15130, B2 => REGISTERS_16_43_port, ZN => n14201);
   U12390 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_43_port, B1 => 
                           n15144, B2 => REGISTERS_9_43_port, ZN => n14200);
   U12391 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_43_port, B1 => 
                           n15032, B2 => REGISTERS_30_43_port, ZN => n14199);
   U12392 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_43_port, B1 => 
                           n15156, B2 => REGISTERS_23_43_port, ZN => n14198);
   U12393 : NAND4_X1 port map( A1 => n14201, A2 => n14200, A3 => n14199, A4 => 
                           n14198, ZN => n14202);
   U12394 : NOR3_X1 port map( A1 => n14204, A2 => n14203, A3 => n14202, ZN => 
                           n14205);
   U12395 : OAI222_X1 port map( A1 => n16071, A2 => n8485, B1 => n15115, B2 => 
                           n14206, C1 => n14354, C2 => n14205, ZN => n8526);
   U12396 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_42_port, B1 => 
                           n14483, B2 => REGISTERS_4_42_port, ZN => n14210);
   U12397 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_42_port, B1 => 
                           n15090, B2 => REGISTERS_3_42_port, ZN => n14209);
   U12398 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_42_port, B1 => 
                           n15119, B2 => REGISTERS_7_42_port, ZN => n14208);
   U12399 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_42_port, B1 => 
                           n15089, B2 => REGISTERS_0_42_port, ZN => n14207);
   U12400 : AND4_X1 port map( A1 => n14210, A2 => n14209, A3 => n14208, A4 => 
                           n14207, ZN => n14227);
   U12401 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_42_port, B1 => 
                           n15144, B2 => REGISTERS_9_42_port, ZN => n14214);
   U12402 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_42_port, B1 => 
                           n15130, B2 => REGISTERS_16_42_port, ZN => n14213);
   U12403 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_42_port, B1 => 
                           n15142, B2 => REGISTERS_14_42_port, ZN => n14212);
   U12404 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_42_port, B1 => 
                           n15152, B2 => REGISTERS_31_42_port, ZN => n14211);
   U12405 : NAND4_X1 port map( A1 => n14214, A2 => n14213, A3 => n14212, A4 => 
                           n14211, ZN => n14225);
   U12406 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_42_port, B1 => 
                           n15128, B2 => REGISTERS_22_42_port, ZN => n14218);
   U12407 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_42_port, B1 => 
                           n15127, B2 => REGISTERS_24_42_port, ZN => n14217);
   U12408 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_42_port, B1 => 
                           n14837, B2 => REGISTERS_28_42_port, ZN => n14216);
   U12409 : AOI22_X1 port map( A1 => n14257, A2 => REGISTERS_18_42_port, B1 => 
                           n15140, B2 => REGISTERS_12_42_port, ZN => n14215);
   U12410 : NAND4_X1 port map( A1 => n14218, A2 => n14217, A3 => n14216, A4 => 
                           n14215, ZN => n14224);
   U12411 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_42_port, B1 => 
                           n15150, B2 => REGISTERS_10_42_port, ZN => n14222);
   U12412 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_42_port, B1 => 
                           n15154, B2 => REGISTERS_21_42_port, ZN => n14221);
   U12413 : AOI22_X1 port map( A1 => n15145, A2 => REGISTERS_8_42_port, B1 => 
                           n15126, B2 => REGISTERS_29_42_port, ZN => n14220);
   U12414 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_42_port, B1 => 
                           n15143, B2 => REGISTERS_27_42_port, ZN => n14219);
   U12415 : NAND4_X1 port map( A1 => n14222, A2 => n14221, A3 => n14220, A4 => 
                           n14219, ZN => n14223);
   U12416 : NOR3_X1 port map( A1 => n14225, A2 => n14224, A3 => n14223, ZN => 
                           n14226);
   U12417 : OAI222_X1 port map( A1 => n16071, A2 => n8484, B1 => n14505, B2 => 
                           n14227, C1 => n14354, C2 => n14226, ZN => n8527);
   U12418 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_41_port, B1 => 
                           n15121, B2 => REGISTERS_3_41_port, ZN => n14231);
   U12419 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_41_port, B1 => 
                           n15119, B2 => REGISTERS_7_41_port, ZN => n14230);
   U12420 : AOI22_X1 port map( A1 => n14781, A2 => REGISTERS_6_41_port, B1 => 
                           n14483, B2 => REGISTERS_4_41_port, ZN => n14229);
   U12421 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_41_port, B1 => 
                           n15089, B2 => REGISTERS_0_41_port, ZN => n14228);
   U12422 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_41_port, B1 => 
                           n15128, B2 => REGISTERS_22_41_port, ZN => n14235);
   U12423 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_41_port, B1 => 
                           n15096, B2 => REGISTERS_28_41_port, ZN => n14234);
   U12424 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_41_port, B1 => 
                           n15154, B2 => REGISTERS_21_41_port, ZN => n14233);
   U12425 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_41_port, B1 => 
                           n15130, B2 => REGISTERS_16_41_port, ZN => n14232);
   U12426 : NAND4_X1 port map( A1 => n14235, A2 => n14234, A3 => n14233, A4 => 
                           n14232, ZN => n14246);
   U12427 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_41_port, B1 => 
                           n15152, B2 => REGISTERS_31_41_port, ZN => n14239);
   U12428 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_41_port, B1 => 
                           n15153, B2 => REGISTERS_20_41_port, ZN => n14238);
   U12429 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_41_port, B1 => 
                           n14979, B2 => REGISTERS_19_41_port, ZN => n14237);
   U12430 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_41_port, B1 => 
                           n15126, B2 => REGISTERS_29_41_port, ZN => n14236);
   U12431 : NAND4_X1 port map( A1 => n14239, A2 => n14238, A3 => n14237, A4 => 
                           n14236, ZN => n14245);
   U12432 : AOI22_X1 port map( A1 => n15142, A2 => REGISTERS_14_41_port, B1 => 
                           n15145, B2 => REGISTERS_8_41_port, ZN => n14243);
   U12433 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_41_port, B1 => 
                           n15144, B2 => REGISTERS_9_41_port, ZN => n14242);
   U12434 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_41_port, B1 => 
                           n15127, B2 => REGISTERS_24_41_port, ZN => n14241);
   U12435 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_41_port, B1 => 
                           n15140, B2 => REGISTERS_12_41_port, ZN => n14240);
   U12436 : NAND4_X1 port map( A1 => n14243, A2 => n14242, A3 => n14241, A4 => 
                           n14240, ZN => n14244);
   U12437 : NOR3_X1 port map( A1 => n14246, A2 => n14245, A3 => n14244, ZN => 
                           n14247);
   U12438 : OAI222_X1 port map( A1 => n16071, A2 => n8483, B1 => n14505, B2 => 
                           n14248, C1 => n14354, C2 => n14247, ZN => n8528);
   U12439 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_40_port, B1 => 
                           n15119, B2 => REGISTERS_7_40_port, ZN => n14252);
   U12440 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_40_port, B1 => 
                           n15089, B2 => REGISTERS_0_40_port, ZN => n14251);
   U12441 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_40_port, B1 => 
                           n14483, B2 => REGISTERS_4_40_port, ZN => n14250);
   U12442 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_40_port, B1 => 
                           n15065, B2 => REGISTERS_1_40_port, ZN => n14249);
   U12443 : AND4_X1 port map( A1 => n14252, A2 => n14251, A3 => n14250, A4 => 
                           n14249, ZN => n14270);
   U12444 : AOI22_X1 port map( A1 => n15126, A2 => REGISTERS_29_40_port, B1 => 
                           n15154, B2 => REGISTERS_21_40_port, ZN => n14256);
   U12445 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_40_port, B1 => 
                           n15151, B2 => REGISTERS_28_40_port, ZN => n14255);
   U12446 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_40_port, B1 => 
                           n15142, B2 => REGISTERS_14_40_port, ZN => n14254);
   U12447 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_40_port, B1 => 
                           n15156, B2 => REGISTERS_23_40_port, ZN => n14253);
   U12448 : NAND4_X1 port map( A1 => n14256, A2 => n14255, A3 => n14254, A4 => 
                           n14253, ZN => n14268);
   U12449 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_40_port, B1 => 
                           n15139, B2 => REGISTERS_19_40_port, ZN => n14261);
   U12450 : AOI22_X1 port map( A1 => n14257, A2 => REGISTERS_18_40_port, B1 => 
                           n15130, B2 => REGISTERS_16_40_port, ZN => n14260);
   U12451 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_40_port, B1 => 
                           n15145, B2 => REGISTERS_8_40_port, ZN => n14259);
   U12452 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_40_port, B1 => 
                           n15150, B2 => REGISTERS_10_40_port, ZN => n14258);
   U12453 : NAND4_X1 port map( A1 => n14261, A2 => n14260, A3 => n14259, A4 => 
                           n14258, ZN => n14267);
   U12454 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_40_port, B1 => 
                           n15127, B2 => REGISTERS_24_40_port, ZN => n14265);
   U12455 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_40_port, B1 => 
                           n15144, B2 => REGISTERS_9_40_port, ZN => n14264);
   U12456 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_40_port, B1 => 
                           n15138, B2 => REGISTERS_11_40_port, ZN => n14263);
   U12457 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_40_port, B1 => 
                           n15128, B2 => REGISTERS_22_40_port, ZN => n14262);
   U12458 : NAND4_X1 port map( A1 => n14265, A2 => n14264, A3 => n14263, A4 => 
                           n14262, ZN => n14266);
   U12459 : NOR3_X1 port map( A1 => n14268, A2 => n14267, A3 => n14266, ZN => 
                           n14269);
   U12460 : OAI222_X1 port map( A1 => n16071, A2 => n8482, B1 => n14505, B2 => 
                           n14270, C1 => n14354, C2 => n14269, ZN => n8529);
   U12461 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_39_port, B1 => 
                           n14483, B2 => REGISTERS_4_39_port, ZN => n14274);
   U12462 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_39_port, B1 => 
                           n15119, B2 => REGISTERS_7_39_port, ZN => n14273);
   U12463 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_39_port, B1 => 
                           n15089, B2 => REGISTERS_0_39_port, ZN => n14272);
   U12464 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_39_port, B1 => 
                           n15043, B2 => REGISTERS_6_39_port, ZN => n14271);
   U12465 : AND4_X1 port map( A1 => n14274, A2 => n14273, A3 => n14272, A4 => 
                           n14271, ZN => n14291);
   U12466 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_39_port, B1 => 
                           n15142, B2 => REGISTERS_14_39_port, ZN => n14278);
   U12467 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_39_port, B1 => 
                           n15156, B2 => REGISTERS_23_39_port, ZN => n14277);
   U12468 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_39_port, B1 => 
                           n15145, B2 => REGISTERS_8_39_port, ZN => n14276);
   U12469 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_39_port, B1 => 
                           n15152, B2 => REGISTERS_31_39_port, ZN => n14275);
   U12470 : NAND4_X1 port map( A1 => n14278, A2 => n14277, A3 => n14276, A4 => 
                           n14275, ZN => n14289);
   U12471 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_39_port, B1 => 
                           n15130, B2 => REGISTERS_16_39_port, ZN => n14282);
   U12472 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_39_port, B1 => 
                           n14944, B2 => REGISTERS_25_39_port, ZN => n14281);
   U12473 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_39_port, B1 => 
                           n15096, B2 => REGISTERS_28_39_port, ZN => n14280);
   U12474 : AOI22_X1 port map( A1 => n15126, A2 => REGISTERS_29_39_port, B1 => 
                           n15128, B2 => REGISTERS_22_39_port, ZN => n14279);
   U12475 : NAND4_X1 port map( A1 => n14282, A2 => n14281, A3 => n14280, A4 => 
                           n14279, ZN => n14288);
   U12476 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_39_port, B1 => 
                           n15138, B2 => REGISTERS_11_39_port, ZN => n14286);
   U12477 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_39_port, B1 => 
                           n15154, B2 => REGISTERS_21_39_port, ZN => n14285);
   U12478 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_39_port, B1 => 
                           n15127, B2 => REGISTERS_24_39_port, ZN => n14284);
   U12479 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_39_port, B1 => 
                           n15144, B2 => REGISTERS_9_39_port, ZN => n14283);
   U12480 : NAND4_X1 port map( A1 => n14286, A2 => n14285, A3 => n14284, A4 => 
                           n14283, ZN => n14287);
   U12481 : NOR3_X1 port map( A1 => n14289, A2 => n14288, A3 => n14287, ZN => 
                           n14290);
   U12482 : OAI222_X1 port map( A1 => n16071, A2 => n8481, B1 => n14505, B2 => 
                           n14291, C1 => n14354, C2 => n14290, ZN => n8530);
   U12483 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_38_port, B1 => 
                           n14483, B2 => REGISTERS_4_38_port, ZN => n14295);
   U12484 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_38_port, B1 => 
                           n15091, B2 => REGISTERS_7_38_port, ZN => n14294);
   U12485 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_38_port, B1 => 
                           n15089, B2 => REGISTERS_0_38_port, ZN => n14293);
   U12486 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_38_port, B1 => 
                           n14781, B2 => REGISTERS_6_38_port, ZN => n14292);
   U12487 : AND4_X1 port map( A1 => n14295, A2 => n14294, A3 => n14293, A4 => 
                           n14292, ZN => n14312);
   U12488 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_38_port, B1 => 
                           n15126, B2 => REGISTERS_29_38_port, ZN => n14299);
   U12489 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_38_port, B1 => 
                           n15145, B2 => REGISTERS_8_38_port, ZN => n14298);
   U12490 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_38_port, B1 => 
                           n15154, B2 => REGISTERS_21_38_port, ZN => n14297);
   U12491 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_38_port, B1 => 
                           n15128, B2 => REGISTERS_22_38_port, ZN => n14296);
   U12492 : NAND4_X1 port map( A1 => n14299, A2 => n14298, A3 => n14297, A4 => 
                           n14296, ZN => n14310);
   U12493 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_38_port, B1 => 
                           n15144, B2 => REGISTERS_9_38_port, ZN => n14303);
   U12494 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_38_port, B1 => 
                           n15140, B2 => REGISTERS_12_38_port, ZN => n14302);
   U12495 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_38_port, B1 => 
                           n15132, B2 => REGISTERS_15_38_port, ZN => n14301);
   U12496 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_38_port, B1 => 
                           n15142, B2 => REGISTERS_14_38_port, ZN => n14300);
   U12497 : NAND4_X1 port map( A1 => n14303, A2 => n14302, A3 => n14301, A4 => 
                           n14300, ZN => n14309);
   U12498 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_38_port, B1 => 
                           n15153, B2 => REGISTERS_20_38_port, ZN => n14307);
   U12499 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_38_port, B1 => 
                           n15150, B2 => REGISTERS_10_38_port, ZN => n14306);
   U12500 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_38_port, B1 => 
                           n15096, B2 => REGISTERS_28_38_port, ZN => n14305);
   U12501 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_38_port, B1 => 
                           n15130, B2 => REGISTERS_16_38_port, ZN => n14304);
   U12502 : NAND4_X1 port map( A1 => n14307, A2 => n14306, A3 => n14305, A4 => 
                           n14304, ZN => n14308);
   U12503 : NOR3_X1 port map( A1 => n14310, A2 => n14309, A3 => n14308, ZN => 
                           n14311);
   U12504 : OAI222_X1 port map( A1 => n16071, A2 => n8480, B1 => n15115, B2 => 
                           n14312, C1 => n14354, C2 => n14311, ZN => n8531);
   U12505 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_37_port, B1 => 
                           n15090, B2 => REGISTERS_3_37_port, ZN => n14316);
   U12506 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_37_port, B1 => 
                           n15089, B2 => REGISTERS_0_37_port, ZN => n14315);
   U12507 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_37_port, B1 => 
                           n15091, B2 => REGISTERS_7_37_port, ZN => n14314);
   U12508 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_37_port, B1 => 
                           n14483, B2 => REGISTERS_4_37_port, ZN => n14313);
   U12509 : AND4_X1 port map( A1 => n14316, A2 => n14315, A3 => n14314, A4 => 
                           n14313, ZN => n14333);
   U12510 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_37_port, B1 => 
                           n15032, B2 => REGISTERS_30_37_port, ZN => n14320);
   U12511 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_37_port, B1 => 
                           n15132, B2 => REGISTERS_15_37_port, ZN => n14319);
   U12512 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_37_port, B1 => 
                           n15144, B2 => REGISTERS_9_37_port, ZN => n14318);
   U12513 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_37_port, B1 => 
                           n15127, B2 => REGISTERS_24_37_port, ZN => n14317);
   U12514 : NAND4_X1 port map( A1 => n14320, A2 => n14319, A3 => n14318, A4 => 
                           n14317, ZN => n14331);
   U12515 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_37_port, B1 => 
                           n15145, B2 => REGISTERS_8_37_port, ZN => n14324);
   U12516 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_37_port, B1 => 
                           n15142, B2 => REGISTERS_14_37_port, ZN => n14323);
   U12517 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_37_port, B1 => 
                           n15154, B2 => REGISTERS_21_37_port, ZN => n14322);
   U12518 : AOI22_X1 port map( A1 => n15126, A2 => REGISTERS_29_37_port, B1 => 
                           n15128, B2 => REGISTERS_22_37_port, ZN => n14321);
   U12519 : NAND4_X1 port map( A1 => n14324, A2 => n14323, A3 => n14322, A4 => 
                           n14321, ZN => n14330);
   U12520 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_37_port, B1 => 
                           n14837, B2 => REGISTERS_28_37_port, ZN => n14328);
   U12521 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_37_port, B1 => 
                           n15150, B2 => REGISTERS_10_37_port, ZN => n14327);
   U12522 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_37_port, B1 => 
                           n15140, B2 => REGISTERS_12_37_port, ZN => n14326);
   U12523 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_37_port, B1 => 
                           n15152, B2 => REGISTERS_31_37_port, ZN => n14325);
   U12524 : NAND4_X1 port map( A1 => n14328, A2 => n14327, A3 => n14326, A4 => 
                           n14325, ZN => n14329);
   U12525 : NOR3_X1 port map( A1 => n14331, A2 => n14330, A3 => n14329, ZN => 
                           n14332);
   U12526 : OAI222_X1 port map( A1 => n16071, A2 => n8479, B1 => n14505, B2 => 
                           n14333, C1 => n14354, C2 => n14332, ZN => n8532);
   U12527 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_36_port, B1 => 
                           n15089, B2 => REGISTERS_0_36_port, ZN => n14337);
   U12528 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_36_port, B1 => 
                           n15091, B2 => REGISTERS_7_36_port, ZN => n14336);
   U12529 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_36_port, B1 => 
                           n15043, B2 => REGISTERS_6_36_port, ZN => n14335);
   U12530 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_36_port, B1 => 
                           n14483, B2 => REGISTERS_4_36_port, ZN => n14334);
   U12531 : AND4_X1 port map( A1 => n14337, A2 => n14336, A3 => n14335, A4 => 
                           n14334, ZN => n14355);
   U12532 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_36_port, B1 => 
                           n15138, B2 => REGISTERS_11_36_port, ZN => n14341);
   U12533 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_36_port, B1 => 
                           n15152, B2 => REGISTERS_31_36_port, ZN => n14340);
   U12534 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_36_port, B1 => 
                           n15032, B2 => REGISTERS_30_36_port, ZN => n14339);
   U12535 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_36_port, B1 => 
                           n15145, B2 => REGISTERS_8_36_port, ZN => n14338);
   U12536 : NAND4_X1 port map( A1 => n14341, A2 => n14340, A3 => n14339, A4 => 
                           n14338, ZN => n14352);
   U12537 : AOI22_X1 port map( A1 => n15144, A2 => REGISTERS_9_36_port, B1 => 
                           n15154, B2 => REGISTERS_21_36_port, ZN => n14345);
   U12538 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_36_port, B1 => 
                           n15127, B2 => REGISTERS_24_36_port, ZN => n14344);
   U12539 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_36_port, B1 => 
                           n15142, B2 => REGISTERS_14_36_port, ZN => n14343);
   U12540 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_36_port, B1 => 
                           n15153, B2 => REGISTERS_20_36_port, ZN => n14342);
   U12541 : NAND4_X1 port map( A1 => n14345, A2 => n14344, A3 => n14343, A4 => 
                           n14342, ZN => n14351);
   U12542 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_36_port, B1 => 
                           n15150, B2 => REGISTERS_10_36_port, ZN => n14349);
   U12543 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_36_port, B1 => 
                           n15151, B2 => REGISTERS_28_36_port, ZN => n14348);
   U12544 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_36_port, B1 => 
                           n15132, B2 => REGISTERS_15_36_port, ZN => n14347);
   U12545 : AOI22_X1 port map( A1 => n15126, A2 => REGISTERS_29_36_port, B1 => 
                           n15128, B2 => REGISTERS_22_36_port, ZN => n14346);
   U12546 : NAND4_X1 port map( A1 => n14349, A2 => n14348, A3 => n14347, A4 => 
                           n14346, ZN => n14350);
   U12547 : NOR3_X1 port map( A1 => n14352, A2 => n14351, A3 => n14350, ZN => 
                           n14353);
   U12548 : OAI222_X1 port map( A1 => n16071, A2 => n8478, B1 => n15115, B2 => 
                           n14355, C1 => n14354, C2 => n14353, ZN => n8533);
   U12549 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_35_port, B1 => 
                           n14781, B2 => REGISTERS_6_35_port, ZN => n14359);
   U12550 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_35_port, B1 => 
                           n14483, B2 => REGISTERS_4_35_port, ZN => n14358);
   U12551 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_35_port, B1 => 
                           n15089, B2 => REGISTERS_0_35_port, ZN => n14357);
   U12552 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_35_port, B1 => 
                           n15091, B2 => REGISTERS_7_35_port, ZN => n14356);
   U12553 : AND4_X1 port map( A1 => n14359, A2 => n14358, A3 => n14357, A4 => 
                           n14356, ZN => n14376);
   U12554 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_35_port, B1 => 
                           n15153, B2 => REGISTERS_20_35_port, ZN => n14363);
   U12555 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_35_port, B1 => 
                           n15130, B2 => REGISTERS_16_35_port, ZN => n14362);
   U12556 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_35_port, B1 => 
                           n15140, B2 => REGISTERS_12_35_port, ZN => n14361);
   U12557 : AOI22_X1 port map( A1 => n15142, A2 => REGISTERS_14_35_port, B1 => 
                           n15150, B2 => REGISTERS_10_35_port, ZN => n14360);
   U12558 : NAND4_X1 port map( A1 => n14363, A2 => n14362, A3 => n14361, A4 => 
                           n14360, ZN => n14374);
   U12559 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_35_port, B1 => 
                           n15144, B2 => REGISTERS_9_35_port, ZN => n14367);
   U12560 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_35_port, B1 => 
                           n15145, B2 => REGISTERS_8_35_port, ZN => n14366);
   U12561 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_35_port, B1 => 
                           n15139, B2 => REGISTERS_19_35_port, ZN => n14365);
   U12562 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_35_port, B1 => 
                           n15096, B2 => REGISTERS_28_35_port, ZN => n14364);
   U12563 : NAND4_X1 port map( A1 => n14367, A2 => n14366, A3 => n14365, A4 => 
                           n14364, ZN => n14373);
   U12564 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_35_port, B1 => 
                           n15154, B2 => REGISTERS_21_35_port, ZN => n14371);
   U12565 : AOI22_X1 port map( A1 => n15126, A2 => REGISTERS_29_35_port, B1 => 
                           n15128, B2 => REGISTERS_22_35_port, ZN => n14370);
   U12566 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_35_port, B1 => 
                           n15155, B2 => REGISTERS_18_35_port, ZN => n14369);
   U12567 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_35_port, B1 => 
                           n15132, B2 => REGISTERS_15_35_port, ZN => n14368);
   U12568 : NAND4_X1 port map( A1 => n14371, A2 => n14370, A3 => n14369, A4 => 
                           n14368, ZN => n14372);
   U12569 : NOR3_X1 port map( A1 => n14374, A2 => n14373, A3 => n14372, ZN => 
                           n14375);
   U12570 : OAI222_X1 port map( A1 => n16071, A2 => n8477, B1 => n14505, B2 => 
                           n14376, C1 => n14354, C2 => n14375, ZN => n8534);
   U12571 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_34_port, B1 => 
                           n14781, B2 => REGISTERS_6_34_port, ZN => n14380);
   U12572 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_34_port, B1 => 
                           n15089, B2 => REGISTERS_0_34_port, ZN => n14379);
   U12573 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_34_port, B1 => 
                           n15091, B2 => REGISTERS_7_34_port, ZN => n14378);
   U12574 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_34_port, B1 => 
                           n14483, B2 => REGISTERS_4_34_port, ZN => n14377);
   U12575 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_34_port, B1 => 
                           n15139, B2 => REGISTERS_19_34_port, ZN => n14384);
   U12576 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_34_port, B1 => 
                           n15126, B2 => REGISTERS_29_34_port, ZN => n14383);
   U12577 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_34_port, B1 => 
                           n14837, B2 => REGISTERS_28_34_port, ZN => n14382);
   U12578 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_34_port, B1 => 
                           n15154, B2 => REGISTERS_21_34_port, ZN => n14381);
   U12579 : NAND4_X1 port map( A1 => n14384, A2 => n14383, A3 => n14382, A4 => 
                           n14381, ZN => n14395);
   U12580 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_34_port, B1 => 
                           n15156, B2 => REGISTERS_23_34_port, ZN => n14388);
   U12581 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_34_port, B1 => 
                           n15153, B2 => REGISTERS_20_34_port, ZN => n14387);
   U12582 : AOI22_X1 port map( A1 => n15145, A2 => REGISTERS_8_34_port, B1 => 
                           n15128, B2 => REGISTERS_22_34_port, ZN => n14386);
   U12583 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_34_port, B1 => 
                           n15152, B2 => REGISTERS_31_34_port, ZN => n14385);
   U12584 : NAND4_X1 port map( A1 => n14388, A2 => n14387, A3 => n14386, A4 => 
                           n14385, ZN => n14394);
   U12585 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_34_port, B1 => 
                           n15144, B2 => REGISTERS_9_34_port, ZN => n14392);
   U12586 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_34_port, B1 => 
                           n15142, B2 => REGISTERS_14_34_port, ZN => n14391);
   U12587 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_34_port, B1 => 
                           n15130, B2 => REGISTERS_16_34_port, ZN => n14390);
   U12588 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_34_port, B1 => 
                           n15138, B2 => REGISTERS_11_34_port, ZN => n14389);
   U12589 : NAND4_X1 port map( A1 => n14392, A2 => n14391, A3 => n14390, A4 => 
                           n14389, ZN => n14393);
   U12590 : NOR3_X1 port map( A1 => n14395, A2 => n14394, A3 => n14393, ZN => 
                           n14396);
   U12591 : OAI222_X1 port map( A1 => n16071, A2 => n8476, B1 => n15115, B2 => 
                           n14397, C1 => n14354, C2 => n14396, ZN => n8535);
   U12592 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_33_port, B1 => 
                           n15043, B2 => REGISTERS_6_33_port, ZN => n14401);
   U12593 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_33_port, B1 => 
                           n15091, B2 => REGISTERS_7_33_port, ZN => n14400);
   U12594 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_33_port, B1 => 
                           n15121, B2 => REGISTERS_3_33_port, ZN => n14399);
   U12595 : AOI22_X1 port map( A1 => n14483, A2 => REGISTERS_4_33_port, B1 => 
                           n15089, B2 => REGISTERS_0_33_port, ZN => n14398);
   U12596 : AND4_X1 port map( A1 => n14401, A2 => n14400, A3 => n14399, A4 => 
                           n14398, ZN => n14418);
   U12597 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_33_port, B1 => 
                           n15154, B2 => REGISTERS_21_33_port, ZN => n14405);
   U12598 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_33_port, B1 => 
                           n15150, B2 => REGISTERS_10_33_port, ZN => n14404);
   U12599 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_33_port, B1 => 
                           n15145, B2 => REGISTERS_8_33_port, ZN => n14403);
   U12600 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_33_port, B1 => 
                           n15128, B2 => REGISTERS_22_33_port, ZN => n14402);
   U12601 : NAND4_X1 port map( A1 => n14405, A2 => n14404, A3 => n14403, A4 => 
                           n14402, ZN => n14416);
   U12602 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_33_port, B1 => 
                           n15151, B2 => REGISTERS_28_33_port, ZN => n14409);
   U12603 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_33_port, B1 => 
                           n15155, B2 => REGISTERS_18_33_port, ZN => n14408);
   U12604 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_33_port, B1 => 
                           n15152, B2 => REGISTERS_31_33_port, ZN => n14407);
   U12605 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_33_port, B1 => 
                           n15032, B2 => REGISTERS_30_33_port, ZN => n14406);
   U12606 : NAND4_X1 port map( A1 => n14409, A2 => n14408, A3 => n14407, A4 => 
                           n14406, ZN => n14415);
   U12607 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_33_port, B1 => 
                           n15156, B2 => REGISTERS_23_33_port, ZN => n14413);
   U12608 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_33_port, B1 => 
                           n15126, B2 => REGISTERS_29_33_port, ZN => n14412);
   U12609 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_33_port, B1 => 
                           n15142, B2 => REGISTERS_14_33_port, ZN => n14411);
   U12610 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_33_port, B1 => 
                           n15144, B2 => REGISTERS_9_33_port, ZN => n14410);
   U12611 : NAND4_X1 port map( A1 => n14413, A2 => n14412, A3 => n14411, A4 => 
                           n14410, ZN => n14414);
   U12612 : NOR3_X1 port map( A1 => n14416, A2 => n14415, A3 => n14414, ZN => 
                           n14417);
   U12613 : OAI222_X1 port map( A1 => n16071, A2 => n8475, B1 => n14505, B2 => 
                           n14418, C1 => n15166, C2 => n14417, ZN => n8536);
   U12614 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_32_port, B1 => 
                           n14483, B2 => REGISTERS_4_32_port, ZN => n14422);
   U12615 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_32_port, B1 => 
                           n15089, B2 => REGISTERS_0_32_port, ZN => n14421);
   U12616 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_32_port, B1 => 
                           n15091, B2 => REGISTERS_7_32_port, ZN => n14420);
   U12617 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_32_port, B1 => 
                           n15043, B2 => REGISTERS_6_32_port, ZN => n14419);
   U12618 : AND4_X1 port map( A1 => n14422, A2 => n14421, A3 => n14420, A4 => 
                           n14419, ZN => n14439);
   U12619 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_32_port, B1 => 
                           n15144, B2 => REGISTERS_9_32_port, ZN => n14426);
   U12620 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_32_port, B1 => 
                           n15126, B2 => REGISTERS_29_32_port, ZN => n14425);
   U12621 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_32_port, B1 => 
                           n15152, B2 => REGISTERS_31_32_port, ZN => n14424);
   U12622 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_32_port, B1 => 
                           n15156, B2 => REGISTERS_23_32_port, ZN => n14423);
   U12623 : NAND4_X1 port map( A1 => n14426, A2 => n14425, A3 => n14424, A4 => 
                           n14423, ZN => n14437);
   U12624 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_32_port, B1 => 
                           n15142, B2 => REGISTERS_14_32_port, ZN => n14430);
   U12625 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_32_port, B1 => 
                           n15138, B2 => REGISTERS_11_32_port, ZN => n14429);
   U12626 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_32_port, B1 => 
                           n15032, B2 => REGISTERS_30_32_port, ZN => n14428);
   U12627 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_32_port, B1 => 
                           n15145, B2 => REGISTERS_8_32_port, ZN => n14427);
   U12628 : NAND4_X1 port map( A1 => n14430, A2 => n14429, A3 => n14428, A4 => 
                           n14427, ZN => n14436);
   U12629 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_32_port, B1 => 
                           n15154, B2 => REGISTERS_21_32_port, ZN => n14434);
   U12630 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_32_port, B1 => 
                           n15096, B2 => REGISTERS_28_32_port, ZN => n14433);
   U12631 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_32_port, B1 => 
                           n15130, B2 => REGISTERS_16_32_port, ZN => n14432);
   U12632 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_32_port, B1 => 
                           n15128, B2 => REGISTERS_22_32_port, ZN => n14431);
   U12633 : NAND4_X1 port map( A1 => n14434, A2 => n14433, A3 => n14432, A4 => 
                           n14431, ZN => n14435);
   U12634 : NOR3_X1 port map( A1 => n14437, A2 => n14436, A3 => n14435, ZN => 
                           n14438);
   U12635 : OAI222_X1 port map( A1 => n16071, A2 => n8474, B1 => n15115, B2 => 
                           n14439, C1 => n14354, C2 => n14438, ZN => n8537);
   U12636 : AOI22_X1 port map( A1 => n15117, A2 => REGISTERS_4_31_port, B1 => 
                           n15091, B2 => REGISTERS_7_31_port, ZN => n14443);
   U12637 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_31_port, B1 => 
                           n14781, B2 => REGISTERS_6_31_port, ZN => n14442);
   U12638 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_31_port, B1 => 
                           n15089, B2 => REGISTERS_0_31_port, ZN => n14441);
   U12639 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_31_port, B1 => 
                           n15065, B2 => REGISTERS_1_31_port, ZN => n14440);
   U12640 : AND4_X1 port map( A1 => n14443, A2 => n14442, A3 => n14441, A4 => 
                           n14440, ZN => n14460);
   U12641 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_31_port, B1 => 
                           n15128, B2 => REGISTERS_22_31_port, ZN => n14447);
   U12642 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_31_port, B1 => 
                           n15142, B2 => REGISTERS_14_31_port, ZN => n14446);
   U12643 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_31_port, B1 => 
                           n15126, B2 => REGISTERS_29_31_port, ZN => n14445);
   U12644 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_31_port, B1 => 
                           n14837, B2 => REGISTERS_28_31_port, ZN => n14444);
   U12645 : NAND4_X1 port map( A1 => n14447, A2 => n14446, A3 => n14445, A4 => 
                           n14444, ZN => n14458);
   U12646 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_31_port, B1 => 
                           n15127, B2 => REGISTERS_24_31_port, ZN => n14451);
   U12647 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_31_port, B1 => 
                           n15152, B2 => REGISTERS_31_31_port, ZN => n14450);
   U12648 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_31_port, B1 => 
                           n15145, B2 => REGISTERS_8_31_port, ZN => n14449);
   U12649 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_31_port, B1 => 
                           n15150, B2 => REGISTERS_10_31_port, ZN => n14448);
   U12650 : NAND4_X1 port map( A1 => n14451, A2 => n14450, A3 => n14449, A4 => 
                           n14448, ZN => n14457);
   U12651 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_31_port, B1 => 
                           n15154, B2 => REGISTERS_21_31_port, ZN => n14455);
   U12652 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_31_port, B1 => 
                           n15132, B2 => REGISTERS_15_31_port, ZN => n14454);
   U12653 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_31_port, B1 => 
                           n15074, B2 => REGISTERS_30_31_port, ZN => n14453);
   U12654 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_31_port, B1 => 
                           n15144, B2 => REGISTERS_9_31_port, ZN => n14452);
   U12655 : NAND4_X1 port map( A1 => n14455, A2 => n14454, A3 => n14453, A4 => 
                           n14452, ZN => n14456);
   U12656 : NOR3_X1 port map( A1 => n14458, A2 => n14457, A3 => n14456, ZN => 
                           n14459);
   U12657 : OAI222_X1 port map( A1 => n16026, A2 => n8473, B1 => n14505, B2 => 
                           n14460, C1 => n14354, C2 => n14459, ZN => n8538);
   U12658 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_30_port, B1 => 
                           n15088, B2 => REGISTERS_5_30_port, ZN => n14465);
   U12659 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_30_port, B1 => 
                           n15121, B2 => REGISTERS_3_30_port, ZN => n14464);
   U12660 : AOI22_X1 port map( A1 => n15117, A2 => REGISTERS_4_30_port, B1 => 
                           n15089, B2 => REGISTERS_0_30_port, ZN => n14463);
   U12661 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_30_port, B1 => 
                           n15119, B2 => REGISTERS_7_30_port, ZN => n14462);
   U12662 : AND4_X1 port map( A1 => n14465, A2 => n14464, A3 => n14463, A4 => 
                           n14462, ZN => n14482);
   U12663 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_30_port, B1 => 
                           n15154, B2 => REGISTERS_21_30_port, ZN => n14469);
   U12664 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_30_port, B1 => 
                           n15126, B2 => REGISTERS_29_30_port, ZN => n14468);
   U12665 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_30_port, B1 => 
                           n14979, B2 => REGISTERS_19_30_port, ZN => n14467);
   U12666 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_30_port, B1 => 
                           n15138, B2 => REGISTERS_11_30_port, ZN => n14466);
   U12667 : NAND4_X1 port map( A1 => n14469, A2 => n14468, A3 => n14467, A4 => 
                           n14466, ZN => n14480);
   U12668 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_30_port, B1 => 
                           n15132, B2 => REGISTERS_15_30_port, ZN => n14473);
   U12669 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_30_port, B1 => 
                           n15127, B2 => REGISTERS_24_30_port, ZN => n14472);
   U12670 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_30_port, B1 => 
                           n15152, B2 => REGISTERS_31_30_port, ZN => n14471);
   U12671 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_30_port, B1 => 
                           n15144, B2 => REGISTERS_9_30_port, ZN => n14470);
   U12672 : NAND4_X1 port map( A1 => n14473, A2 => n14472, A3 => n14471, A4 => 
                           n14470, ZN => n14479);
   U12673 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_30_port, B1 => 
                           n15142, B2 => REGISTERS_14_30_port, ZN => n14477);
   U12674 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_30_port, B1 => 
                           n15150, B2 => REGISTERS_10_30_port, ZN => n14476);
   U12675 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_30_port, B1 => 
                           n15128, B2 => REGISTERS_22_30_port, ZN => n14475);
   U12676 : AOI22_X1 port map( A1 => n15151, A2 => REGISTERS_28_30_port, B1 => 
                           n15145, B2 => REGISTERS_8_30_port, ZN => n14474);
   U12677 : NAND4_X1 port map( A1 => n14477, A2 => n14476, A3 => n14475, A4 => 
                           n14474, ZN => n14478);
   U12678 : NOR3_X1 port map( A1 => n14480, A2 => n14479, A3 => n14478, ZN => 
                           n14481);
   U12679 : OAI222_X1 port map( A1 => n16071, A2 => n8472, B1 => n15115, B2 => 
                           n14482, C1 => n15166, C2 => n14481, ZN => n8539);
   U12680 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_29_port, B1 => 
                           n15089, B2 => REGISTERS_0_29_port, ZN => n14487);
   U12681 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_29_port, B1 => 
                           n15119, B2 => REGISTERS_7_29_port, ZN => n14486);
   U12682 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_29_port, B1 => 
                           n14781, B2 => REGISTERS_6_29_port, ZN => n14485);
   U12683 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_29_port, B1 => 
                           n14483, B2 => REGISTERS_4_29_port, ZN => n14484);
   U12684 : AND4_X1 port map( A1 => n14487, A2 => n14486, A3 => n14485, A4 => 
                           n14484, ZN => n14504);
   U12685 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_29_port, B1 => 
                           n15156, B2 => REGISTERS_23_29_port, ZN => n14491);
   U12686 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_29_port, B1 => 
                           n15132, B2 => REGISTERS_15_29_port, ZN => n14490);
   U12687 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_29_port, B1 => 
                           n15152, B2 => REGISTERS_31_29_port, ZN => n14489);
   U12688 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_29_port, B1 => 
                           n15128, B2 => REGISTERS_22_29_port, ZN => n14488);
   U12689 : NAND4_X1 port map( A1 => n14491, A2 => n14490, A3 => n14489, A4 => 
                           n14488, ZN => n14502);
   U12690 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_29_port, B1 => 
                           n15130, B2 => REGISTERS_16_29_port, ZN => n14495);
   U12691 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_29_port, B1 => 
                           n15154, B2 => REGISTERS_21_29_port, ZN => n14494);
   U12692 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_29_port, B1 => 
                           n15150, B2 => REGISTERS_10_29_port, ZN => n14493);
   U12693 : AOI22_X1 port map( A1 => n15145, A2 => REGISTERS_8_29_port, B1 => 
                           n15144, B2 => REGISTERS_9_29_port, ZN => n14492);
   U12694 : NAND4_X1 port map( A1 => n14495, A2 => n14494, A3 => n14493, A4 => 
                           n14492, ZN => n14501);
   U12695 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_29_port, B1 => 
                           n15142, B2 => REGISTERS_14_29_port, ZN => n14499);
   U12696 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_29_port, B1 => 
                           n15127, B2 => REGISTERS_24_29_port, ZN => n14498);
   U12697 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_29_port, B1 => 
                           n15151, B2 => REGISTERS_28_29_port, ZN => n14497);
   U12698 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_29_port, B1 => 
                           n15126, B2 => REGISTERS_29_29_port, ZN => n14496);
   U12699 : NAND4_X1 port map( A1 => n14499, A2 => n14498, A3 => n14497, A4 => 
                           n14496, ZN => n14500);
   U12700 : NOR3_X1 port map( A1 => n14502, A2 => n14501, A3 => n14500, ZN => 
                           n14503);
   U12701 : OAI222_X1 port map( A1 => n16026, A2 => n8471, B1 => n14505, B2 => 
                           n14504, C1 => n15166, C2 => n14503, ZN => n8540);
   U12702 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_28_port, B1 => 
                           n14781, B2 => REGISTERS_6_28_port, ZN => n14510);
   U12703 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_28_port, B1 => 
                           n15089, B2 => REGISTERS_0_28_port, ZN => n14509);
   U12704 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_28_port, B1 => 
                           n15119, B2 => REGISTERS_7_28_port, ZN => n14508);
   U12705 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_28_port, B1 => 
                           n14483, B2 => REGISTERS_4_28_port, ZN => n14507);
   U12706 : AND4_X1 port map( A1 => n14510, A2 => n14509, A3 => n14508, A4 => 
                           n14507, ZN => n14527);
   U12707 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_28_port, B1 => 
                           n15133, B2 => REGISTERS_30_28_port, ZN => n14514);
   U12708 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_28_port, B1 => 
                           n15127, B2 => REGISTERS_24_28_port, ZN => n14513);
   U12709 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_28_port, B1 => 
                           n15142, B2 => REGISTERS_14_28_port, ZN => n14512);
   U12710 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_28_port, B1 => 
                           n15138, B2 => REGISTERS_11_28_port, ZN => n14511);
   U12711 : NAND4_X1 port map( A1 => n14514, A2 => n14513, A3 => n14512, A4 => 
                           n14511, ZN => n14525);
   U12712 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_28_port, B1 => 
                           n15145, B2 => REGISTERS_8_28_port, ZN => n14518);
   U12713 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_28_port, B1 => 
                           n15152, B2 => REGISTERS_31_28_port, ZN => n14517);
   U12714 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_28_port, B1 => 
                           n15154, B2 => REGISTERS_21_28_port, ZN => n14516);
   U12715 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_28_port, B1 => 
                           n15126, B2 => REGISTERS_29_28_port, ZN => n14515);
   U12716 : NAND4_X1 port map( A1 => n14518, A2 => n14517, A3 => n14516, A4 => 
                           n14515, ZN => n14524);
   U12717 : AOI22_X1 port map( A1 => n15096, A2 => REGISTERS_28_28_port, B1 => 
                           n15144, B2 => REGISTERS_9_28_port, ZN => n14522);
   U12718 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_28_port, B1 => 
                           n15128, B2 => REGISTERS_22_28_port, ZN => n14521);
   U12719 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_28_port, B1 => 
                           n15150, B2 => REGISTERS_10_28_port, ZN => n14520);
   U12720 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_28_port, B1 => 
                           n15153, B2 => REGISTERS_20_28_port, ZN => n14519);
   U12721 : NAND4_X1 port map( A1 => n14522, A2 => n14521, A3 => n14520, A4 => 
                           n14519, ZN => n14523);
   U12722 : NOR3_X1 port map( A1 => n14525, A2 => n14524, A3 => n14523, ZN => 
                           n14526);
   U12723 : OAI222_X1 port map( A1 => n16071, A2 => n8470, B1 => n15115, B2 => 
                           n14527, C1 => n14354, C2 => n14526, ZN => n8541);
   U12724 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_27_port, B1 => 
                           n14781, B2 => REGISTERS_6_27_port, ZN => n14531);
   U12725 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_27_port, B1 => 
                           n15119, B2 => REGISTERS_7_27_port, ZN => n14530);
   U12726 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_27_port, B1 => 
                           n15116, B2 => REGISTERS_0_27_port, ZN => n14529);
   U12727 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_27_port, B1 => 
                           n14483, B2 => REGISTERS_4_27_port, ZN => n14528);
   U12728 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_27_port, B1 => 
                           n15128, B2 => REGISTERS_22_27_port, ZN => n14535);
   U12729 : AOI22_X1 port map( A1 => n15145, A2 => REGISTERS_8_27_port, B1 => 
                           n15126, B2 => REGISTERS_29_27_port, ZN => n14534);
   U12730 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_27_port, B1 => 
                           n15138, B2 => REGISTERS_11_27_port, ZN => n14533);
   U12731 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_27_port, B1 => 
                           n15153, B2 => REGISTERS_20_27_port, ZN => n14532);
   U12732 : NAND4_X1 port map( A1 => n14535, A2 => n14534, A3 => n14533, A4 => 
                           n14532, ZN => n14546);
   U12733 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_27_port, B1 => 
                           n15157, B2 => REGISTERS_13_27_port, ZN => n14539);
   U12734 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_27_port, B1 => 
                           n15142, B2 => REGISTERS_14_27_port, ZN => n14538);
   U12735 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_27_port, B1 => 
                           n15096, B2 => REGISTERS_28_27_port, ZN => n14537);
   U12736 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_27_port, B1 => 
                           n15150, B2 => REGISTERS_10_27_port, ZN => n14536);
   U12737 : NAND4_X1 port map( A1 => n14539, A2 => n14538, A3 => n14537, A4 => 
                           n14536, ZN => n14545);
   U12738 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_27_port, B1 => 
                           n15132, B2 => REGISTERS_15_27_port, ZN => n14543);
   U12739 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_27_port, B1 => 
                           n15152, B2 => REGISTERS_31_27_port, ZN => n14542);
   U12740 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_27_port, B1 => 
                           n15130, B2 => REGISTERS_16_27_port, ZN => n14541);
   U12741 : AOI22_X1 port map( A1 => n15144, A2 => REGISTERS_9_27_port, B1 => 
                           n15154, B2 => REGISTERS_21_27_port, ZN => n14540);
   U12742 : NAND4_X1 port map( A1 => n14543, A2 => n14542, A3 => n14541, A4 => 
                           n14540, ZN => n14544);
   U12743 : NOR3_X1 port map( A1 => n14546, A2 => n14545, A3 => n14544, ZN => 
                           n14547);
   U12744 : OAI222_X1 port map( A1 => n14910, A2 => n8469, B1 => n15115, B2 => 
                           n14548, C1 => n15166, C2 => n14547, ZN => n8542);
   U12745 : AOI22_X1 port map( A1 => n14483, A2 => REGISTERS_4_26_port, B1 => 
                           n15116, B2 => REGISTERS_0_26_port, ZN => n14552);
   U12746 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_26_port, B1 => 
                           n15121, B2 => REGISTERS_3_26_port, ZN => n14551);
   U12747 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_26_port, B1 => 
                           n14781, B2 => REGISTERS_6_26_port, ZN => n14550);
   U12748 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_26_port, B1 => 
                           n15119, B2 => REGISTERS_7_26_port, ZN => n14549);
   U12749 : AND4_X1 port map( A1 => n14552, A2 => n14551, A3 => n14550, A4 => 
                           n14549, ZN => n14569);
   U12750 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_26_port, B1 => 
                           n15129, B2 => REGISTERS_17_26_port, ZN => n14556);
   U12751 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_26_port, B1 => 
                           n15151, B2 => REGISTERS_28_26_port, ZN => n14555);
   U12752 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_26_port, B1 => 
                           n15138, B2 => REGISTERS_11_26_port, ZN => n14554);
   U12753 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_26_port, B1 => 
                           n15133, B2 => REGISTERS_30_26_port, ZN => n14553);
   U12754 : NAND4_X1 port map( A1 => n14556, A2 => n14555, A3 => n14554, A4 => 
                           n14553, ZN => n14567);
   U12755 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_26_port, B1 => 
                           n15152, B2 => REGISTERS_31_26_port, ZN => n14560);
   U12756 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_26_port, B1 => 
                           n15150, B2 => REGISTERS_10_26_port, ZN => n14559);
   U12757 : AOI22_X1 port map( A1 => n15142, A2 => REGISTERS_14_26_port, B1 => 
                           n15128, B2 => REGISTERS_22_26_port, ZN => n14558);
   U12758 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_26_port, B1 => 
                           n15154, B2 => REGISTERS_21_26_port, ZN => n14557);
   U12759 : NAND4_X1 port map( A1 => n14560, A2 => n14559, A3 => n14558, A4 => 
                           n14557, ZN => n14566);
   U12760 : AOI22_X1 port map( A1 => n15145, A2 => REGISTERS_8_26_port, B1 => 
                           n15126, B2 => REGISTERS_29_26_port, ZN => n14564);
   U12761 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_26_port, B1 => 
                           n15156, B2 => REGISTERS_23_26_port, ZN => n14563);
   U12762 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_26_port, B1 => 
                           n15127, B2 => REGISTERS_24_26_port, ZN => n14562);
   U12763 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_26_port, B1 => 
                           n15144, B2 => REGISTERS_9_26_port, ZN => n14561);
   U12764 : NAND4_X1 port map( A1 => n14564, A2 => n14563, A3 => n14562, A4 => 
                           n14561, ZN => n14565);
   U12765 : NOR3_X1 port map( A1 => n14567, A2 => n14566, A3 => n14565, ZN => 
                           n14568);
   U12766 : OAI222_X1 port map( A1 => n16071, A2 => n8468, B1 => n14505, B2 => 
                           n14569, C1 => n14354, C2 => n14568, ZN => n8543);
   U12767 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_25_port, B1 => 
                           n15088, B2 => REGISTERS_5_25_port, ZN => n14573);
   U12768 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_25_port, B1 => 
                           n15121, B2 => REGISTERS_3_25_port, ZN => n14572);
   U12769 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_25_port, B1 => 
                           n15119, B2 => REGISTERS_7_25_port, ZN => n14571);
   U12770 : AOI22_X1 port map( A1 => n15117, A2 => REGISTERS_4_25_port, B1 => 
                           n15116, B2 => REGISTERS_0_25_port, ZN => n14570);
   U12771 : AND4_X1 port map( A1 => n14573, A2 => n14572, A3 => n14571, A4 => 
                           n14570, ZN => n14590);
   U12772 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_25_port, B1 => 
                           n15128, B2 => REGISTERS_22_25_port, ZN => n14577);
   U12773 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_25_port, B1 => 
                           n15157, B2 => REGISTERS_13_25_port, ZN => n14576);
   U12774 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_25_port, B1 => 
                           n15151, B2 => REGISTERS_28_25_port, ZN => n14575);
   U12775 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_25_port, B1 => 
                           n15144, B2 => REGISTERS_9_25_port, ZN => n14574);
   U12776 : NAND4_X1 port map( A1 => n14577, A2 => n14576, A3 => n14575, A4 => 
                           n14574, ZN => n14588);
   U12777 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_25_port, B1 => 
                           n15156, B2 => REGISTERS_23_25_port, ZN => n14581);
   U12778 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_25_port, B1 => 
                           n15153, B2 => REGISTERS_20_25_port, ZN => n14580);
   U12779 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_25_port, B1 => 
                           n15132, B2 => REGISTERS_15_25_port, ZN => n14579);
   U12780 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_25_port, B1 => 
                           n15126, B2 => REGISTERS_29_25_port, ZN => n14578);
   U12781 : NAND4_X1 port map( A1 => n14581, A2 => n14580, A3 => n14579, A4 => 
                           n14578, ZN => n14587);
   U12782 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_25_port, B1 => 
                           n15154, B2 => REGISTERS_21_25_port, ZN => n14585);
   U12783 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_25_port, B1 => 
                           n15145, B2 => REGISTERS_8_25_port, ZN => n14584);
   U12784 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_25_port, B1 => 
                           n15142, B2 => REGISTERS_14_25_port, ZN => n14583);
   U12785 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_25_port, B1 => 
                           n15152, B2 => REGISTERS_31_25_port, ZN => n14582);
   U12786 : NAND4_X1 port map( A1 => n14585, A2 => n14584, A3 => n14583, A4 => 
                           n14582, ZN => n14586);
   U12787 : NOR3_X1 port map( A1 => n14588, A2 => n14587, A3 => n14586, ZN => 
                           n14589);
   U12788 : OAI222_X1 port map( A1 => n16026, A2 => n8467, B1 => n15115, B2 => 
                           n14590, C1 => n15166, C2 => n14589, ZN => n8544);
   U12789 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_24_port, B1 => 
                           n14781, B2 => REGISTERS_6_24_port, ZN => n14594);
   U12790 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_24_port, B1 => 
                           n15116, B2 => REGISTERS_0_24_port, ZN => n14593);
   U12791 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_24_port, B1 => 
                           n15117, B2 => REGISTERS_4_24_port, ZN => n14592);
   U12792 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_24_port, B1 => 
                           n15119, B2 => REGISTERS_7_24_port, ZN => n14591);
   U12793 : AND4_X1 port map( A1 => n14594, A2 => n14593, A3 => n14592, A4 => 
                           n14591, ZN => n14611);
   U12794 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_24_port, B1 => 
                           n15129, B2 => REGISTERS_17_24_port, ZN => n14598);
   U12795 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_24_port, B1 => 
                           n15130, B2 => REGISTERS_16_24_port, ZN => n14597);
   U12796 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_24_port, B1 => 
                           n15150, B2 => REGISTERS_10_24_port, ZN => n14596);
   U12797 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_24_port, B1 => 
                           n15096, B2 => REGISTERS_28_24_port, ZN => n14595);
   U12798 : NAND4_X1 port map( A1 => n14598, A2 => n14597, A3 => n14596, A4 => 
                           n14595, ZN => n14609);
   U12799 : AOI22_X1 port map( A1 => n15145, A2 => REGISTERS_8_24_port, B1 => 
                           n15144, B2 => REGISTERS_9_24_port, ZN => n14602);
   U12800 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_24_port, B1 => 
                           n15140, B2 => REGISTERS_12_24_port, ZN => n14601);
   U12801 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_24_port, B1 => 
                           n15154, B2 => REGISTERS_21_24_port, ZN => n14600);
   U12802 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_24_port, B1 => 
                           n15156, B2 => REGISTERS_23_24_port, ZN => n14599);
   U12803 : NAND4_X1 port map( A1 => n14602, A2 => n14601, A3 => n14600, A4 => 
                           n14599, ZN => n14608);
   U12804 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_24_port, B1 => 
                           n15133, B2 => REGISTERS_30_24_port, ZN => n14606);
   U12805 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_24_port, B1 => 
                           n15126, B2 => REGISTERS_29_24_port, ZN => n14605);
   U12806 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_24_port, B1 => 
                           n15153, B2 => REGISTERS_20_24_port, ZN => n14604);
   U12807 : AOI22_X1 port map( A1 => n15142, A2 => REGISTERS_14_24_port, B1 => 
                           n15128, B2 => REGISTERS_22_24_port, ZN => n14603);
   U12808 : NAND4_X1 port map( A1 => n14606, A2 => n14605, A3 => n14604, A4 => 
                           n14603, ZN => n14607);
   U12809 : NOR3_X1 port map( A1 => n14609, A2 => n14608, A3 => n14607, ZN => 
                           n14610);
   U12810 : OAI222_X1 port map( A1 => n14910, A2 => n8466, B1 => n14505, B2 => 
                           n14611, C1 => n14354, C2 => n14610, ZN => n8545);
   U12811 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_23_port, B1 => 
                           n15117, B2 => REGISTERS_4_23_port, ZN => n14615);
   U12812 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_23_port, B1 => 
                           n15119, B2 => REGISTERS_7_23_port, ZN => n14614);
   U12813 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_23_port, B1 => 
                           n15116, B2 => REGISTERS_0_23_port, ZN => n14613);
   U12814 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_23_port, B1 => 
                           n15088, B2 => REGISTERS_5_23_port, ZN => n14612);
   U12815 : AND4_X1 port map( A1 => n14615, A2 => n14614, A3 => n14613, A4 => 
                           n14612, ZN => n14632);
   U12816 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_23_port, B1 => 
                           n15141, B2 => REGISTERS_25_23_port, ZN => n14619);
   U12817 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_23_port, B1 => 
                           n15145, B2 => REGISTERS_8_23_port, ZN => n14618);
   U12818 : AOI22_X1 port map( A1 => n15144, A2 => REGISTERS_9_23_port, B1 => 
                           n15128, B2 => REGISTERS_22_23_port, ZN => n14617);
   U12819 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_23_port, B1 => 
                           n15126, B2 => REGISTERS_29_23_port, ZN => n14616);
   U12820 : NAND4_X1 port map( A1 => n14619, A2 => n14618, A3 => n14617, A4 => 
                           n14616, ZN => n14630);
   U12821 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_23_port, B1 => 
                           n15127, B2 => REGISTERS_24_23_port, ZN => n14623);
   U12822 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_23_port, B1 => 
                           n15151, B2 => REGISTERS_28_23_port, ZN => n14622);
   U12823 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_23_port, B1 => 
                           n15156, B2 => REGISTERS_23_23_port, ZN => n14621);
   U12824 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_23_port, B1 => 
                           n15154, B2 => REGISTERS_21_23_port, ZN => n14620);
   U12825 : NAND4_X1 port map( A1 => n14623, A2 => n14622, A3 => n14621, A4 => 
                           n14620, ZN => n14629);
   U12826 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_23_port, B1 => 
                           n15152, B2 => REGISTERS_31_23_port, ZN => n14627);
   U12827 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_23_port, B1 => 
                           n15150, B2 => REGISTERS_10_23_port, ZN => n14626);
   U12828 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_23_port, B1 => 
                           n15132, B2 => REGISTERS_15_23_port, ZN => n14625);
   U12829 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_23_port, B1 => 
                           n15142, B2 => REGISTERS_14_23_port, ZN => n14624);
   U12830 : NAND4_X1 port map( A1 => n14627, A2 => n14626, A3 => n14625, A4 => 
                           n14624, ZN => n14628);
   U12831 : NOR3_X1 port map( A1 => n14630, A2 => n14629, A3 => n14628, ZN => 
                           n14631);
   U12832 : OAI222_X1 port map( A1 => n14910, A2 => n8465, B1 => n15115, B2 => 
                           n14632, C1 => n14354, C2 => n14631, ZN => n8546);
   U12833 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_22_port, B1 => 
                           n15121, B2 => REGISTERS_3_22_port, ZN => n14636);
   U12834 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_22_port, B1 => 
                           n15119, B2 => REGISTERS_7_22_port, ZN => n14635);
   U12835 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_22_port, B1 => 
                           n15116, B2 => REGISTERS_0_22_port, ZN => n14634);
   U12836 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_22_port, B1 => 
                           n15117, B2 => REGISTERS_4_22_port, ZN => n14633);
   U12837 : AND4_X1 port map( A1 => n14636, A2 => n14635, A3 => n14634, A4 => 
                           n14633, ZN => n14653);
   U12838 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_22_port, B1 => 
                           n15126, B2 => REGISTERS_29_22_port, ZN => n14640);
   U12839 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_22_port, B1 => 
                           n15133, B2 => REGISTERS_30_22_port, ZN => n14639);
   U12840 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_22_port, B1 => 
                           n15145, B2 => REGISTERS_8_22_port, ZN => n14638);
   U12841 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_22_port, B1 => 
                           n15140, B2 => REGISTERS_12_22_port, ZN => n14637);
   U12842 : NAND4_X1 port map( A1 => n14640, A2 => n14639, A3 => n14638, A4 => 
                           n14637, ZN => n14651);
   U12843 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_22_port, B1 => 
                           n15127, B2 => REGISTERS_24_22_port, ZN => n14644);
   U12844 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_22_port, B1 => 
                           n15139, B2 => REGISTERS_19_22_port, ZN => n14643);
   U12845 : AOI22_X1 port map( A1 => n15128, A2 => REGISTERS_22_22_port, B1 => 
                           n15154, B2 => REGISTERS_21_22_port, ZN => n14642);
   U12846 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_22_port, B1 => 
                           n15144, B2 => REGISTERS_9_22_port, ZN => n14641);
   U12847 : NAND4_X1 port map( A1 => n14644, A2 => n14643, A3 => n14642, A4 => 
                           n14641, ZN => n14650);
   U12848 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_22_port, B1 => 
                           n15142, B2 => REGISTERS_14_22_port, ZN => n14648);
   U12849 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_22_port, B1 => 
                           n15152, B2 => REGISTERS_31_22_port, ZN => n14647);
   U12850 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_22_port, B1 => 
                           n15153, B2 => REGISTERS_20_22_port, ZN => n14646);
   U12851 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_22_port, B1 => 
                           n14837, B2 => REGISTERS_28_22_port, ZN => n14645);
   U12852 : NAND4_X1 port map( A1 => n14648, A2 => n14647, A3 => n14646, A4 => 
                           n14645, ZN => n14649);
   U12853 : NOR3_X1 port map( A1 => n14651, A2 => n14650, A3 => n14649, ZN => 
                           n14652);
   U12854 : OAI222_X1 port map( A1 => n16071, A2 => n8464, B1 => n14505, B2 => 
                           n14653, C1 => n14354, C2 => n14652, ZN => n8547);
   U12855 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_21_port, B1 => 
                           n15121, B2 => REGISTERS_3_21_port, ZN => n14657);
   U12856 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_21_port, B1 => 
                           n15116, B2 => REGISTERS_0_21_port, ZN => n14656);
   U12857 : AOI22_X1 port map( A1 => n14483, A2 => REGISTERS_4_21_port, B1 => 
                           n15119, B2 => REGISTERS_7_21_port, ZN => n14655);
   U12858 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_21_port, B1 => 
                           n15065, B2 => REGISTERS_1_21_port, ZN => n14654);
   U12859 : AND4_X1 port map( A1 => n14657, A2 => n14656, A3 => n14655, A4 => 
                           n14654, ZN => n14674);
   U12860 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_21_port, B1 => 
                           n15140, B2 => REGISTERS_12_21_port, ZN => n14661);
   U12861 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_21_port, B1 => 
                           n15143, B2 => REGISTERS_27_21_port, ZN => n14660);
   U12862 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_21_port, B1 => 
                           n15127, B2 => REGISTERS_24_21_port, ZN => n14659);
   U12863 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_21_port, B1 => 
                           n15128, B2 => REGISTERS_22_21_port, ZN => n14658);
   U12864 : NAND4_X1 port map( A1 => n14661, A2 => n14660, A3 => n14659, A4 => 
                           n14658, ZN => n14672);
   U12865 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_21_port, B1 => 
                           n15145, B2 => REGISTERS_8_21_port, ZN => n14665);
   U12866 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_21_port, B1 => 
                           n15153, B2 => REGISTERS_20_21_port, ZN => n14664);
   U12867 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_21_port, B1 => 
                           n15096, B2 => REGISTERS_28_21_port, ZN => n14663);
   U12868 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_21_port, B1 => 
                           n15142, B2 => REGISTERS_14_21_port, ZN => n14662);
   U12869 : NAND4_X1 port map( A1 => n14665, A2 => n14664, A3 => n14663, A4 => 
                           n14662, ZN => n14671);
   U12870 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_21_port, B1 => 
                           n15126, B2 => REGISTERS_29_21_port, ZN => n14669);
   U12871 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_21_port, B1 => 
                           n15155, B2 => REGISTERS_18_21_port, ZN => n14668);
   U12872 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_21_port, B1 => 
                           n15154, B2 => REGISTERS_21_21_port, ZN => n14667);
   U12873 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_21_port, B1 => 
                           n15144, B2 => REGISTERS_9_21_port, ZN => n14666);
   U12874 : NAND4_X1 port map( A1 => n14669, A2 => n14668, A3 => n14667, A4 => 
                           n14666, ZN => n14670);
   U12875 : NOR3_X1 port map( A1 => n14672, A2 => n14671, A3 => n14670, ZN => 
                           n14673);
   U12876 : OAI222_X1 port map( A1 => n16026, A2 => n8463, B1 => n15115, B2 => 
                           n14674, C1 => n14354, C2 => n14673, ZN => n8548);
   U12877 : AOI22_X1 port map( A1 => n15117, A2 => REGISTERS_4_20_port, B1 => 
                           n15119, B2 => REGISTERS_7_20_port, ZN => n14678);
   U12878 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_20_port, B1 => 
                           n15065, B2 => REGISTERS_1_20_port, ZN => n14677);
   U12879 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_20_port, B1 => 
                           n15121, B2 => REGISTERS_3_20_port, ZN => n14676);
   U12880 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_20_port, B1 => 
                           n15116, B2 => REGISTERS_0_20_port, ZN => n14675);
   U12881 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_20_port, B1 => 
                           n15153, B2 => REGISTERS_20_20_port, ZN => n14682);
   U12882 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_20_port, B1 => 
                           n15143, B2 => REGISTERS_27_20_port, ZN => n14681);
   U12883 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_20_port, B1 => 
                           n15150, B2 => REGISTERS_10_20_port, ZN => n14680);
   U12884 : AOI22_X1 port map( A1 => n15096, A2 => REGISTERS_28_20_port, B1 => 
                           n15128, B2 => REGISTERS_22_20_port, ZN => n14679);
   U12885 : NAND4_X1 port map( A1 => n14682, A2 => n14681, A3 => n14680, A4 => 
                           n14679, ZN => n14693);
   U12886 : AOI22_X1 port map( A1 => n15142, A2 => REGISTERS_14_20_port, B1 => 
                           n15126, B2 => REGISTERS_29_20_port, ZN => n14686);
   U12887 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_20_port, B1 => 
                           n15138, B2 => REGISTERS_11_20_port, ZN => n14685);
   U12888 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_20_port, B1 => 
                           n15154, B2 => REGISTERS_21_20_port, ZN => n14684);
   U12889 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_20_port, B1 => 
                           n15144, B2 => REGISTERS_9_20_port, ZN => n14683);
   U12890 : NAND4_X1 port map( A1 => n14686, A2 => n14685, A3 => n14684, A4 => 
                           n14683, ZN => n14692);
   U12891 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_20_port, B1 => 
                           n15152, B2 => REGISTERS_31_20_port, ZN => n14690);
   U12892 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_20_port, B1 => 
                           n15140, B2 => REGISTERS_12_20_port, ZN => n14689);
   U12893 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_20_port, B1 => 
                           n15145, B2 => REGISTERS_8_20_port, ZN => n14688);
   U12894 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_20_port, B1 => 
                           n15132, B2 => REGISTERS_15_20_port, ZN => n14687);
   U12895 : NAND4_X1 port map( A1 => n14690, A2 => n14689, A3 => n14688, A4 => 
                           n14687, ZN => n14691);
   U12896 : NOR3_X1 port map( A1 => n14693, A2 => n14692, A3 => n14691, ZN => 
                           n14694);
   U12897 : OAI222_X1 port map( A1 => n14910, A2 => n8462, B1 => n14505, B2 => 
                           n14695, C1 => n14354, C2 => n14694, ZN => n8549);
   U12898 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_19_port, B1 => 
                           n15117, B2 => REGISTERS_4_19_port, ZN => n14699);
   U12899 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_19_port, B1 => 
                           n15116, B2 => REGISTERS_0_19_port, ZN => n14698);
   U12900 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_19_port, B1 => 
                           n15119, B2 => REGISTERS_7_19_port, ZN => n14697);
   U12901 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_19_port, B1 => 
                           n14781, B2 => REGISTERS_6_19_port, ZN => n14696);
   U12902 : AND4_X1 port map( A1 => n14699, A2 => n14698, A3 => n14697, A4 => 
                           n14696, ZN => n14716);
   U12903 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_19_port, B1 => 
                           n15127, B2 => REGISTERS_24_19_port, ZN => n14703);
   U12904 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_19_port, B1 => 
                           n15142, B2 => REGISTERS_14_19_port, ZN => n14702);
   U12905 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_19_port, B1 => 
                           n15138, B2 => REGISTERS_11_19_port, ZN => n14701);
   U12906 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_19_port, B1 => 
                           n15140, B2 => REGISTERS_12_19_port, ZN => n14700);
   U12907 : NAND4_X1 port map( A1 => n14703, A2 => n14702, A3 => n14701, A4 => 
                           n14700, ZN => n14714);
   U12908 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_19_port, B1 => 
                           n14944, B2 => REGISTERS_25_19_port, ZN => n14707);
   U12909 : AOI22_X1 port map( A1 => n15151, A2 => REGISTERS_28_19_port, B1 => 
                           n15126, B2 => REGISTERS_29_19_port, ZN => n14706);
   U12910 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_19_port, B1 => 
                           n15152, B2 => REGISTERS_31_19_port, ZN => n14705);
   U12911 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_19_port, B1 => 
                           n15145, B2 => REGISTERS_8_19_port, ZN => n14704);
   U12912 : NAND4_X1 port map( A1 => n14707, A2 => n14706, A3 => n14705, A4 => 
                           n14704, ZN => n14713);
   U12913 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_19_port, B1 => 
                           n15150, B2 => REGISTERS_10_19_port, ZN => n14711);
   U12914 : AOI22_X1 port map( A1 => n15128, A2 => REGISTERS_22_19_port, B1 => 
                           n15154, B2 => REGISTERS_21_19_port, ZN => n14710);
   U12915 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_19_port, B1 => 
                           n15144, B2 => REGISTERS_9_19_port, ZN => n14709);
   U12916 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_19_port, B1 => 
                           n15130, B2 => REGISTERS_16_19_port, ZN => n14708);
   U12917 : NAND4_X1 port map( A1 => n14711, A2 => n14710, A3 => n14709, A4 => 
                           n14708, ZN => n14712);
   U12918 : NOR3_X1 port map( A1 => n14714, A2 => n14713, A3 => n14712, ZN => 
                           n14715);
   U12919 : OAI222_X1 port map( A1 => n14910, A2 => n8461, B1 => n15115, B2 => 
                           n14716, C1 => n15166, C2 => n14715, ZN => n8550);
   U12920 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_18_port, B1 => 
                           n15116, B2 => REGISTERS_0_18_port, ZN => n14720);
   U12921 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_18_port, B1 => 
                           n14781, B2 => REGISTERS_6_18_port, ZN => n14719);
   U12922 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_18_port, B1 => 
                           n14483, B2 => REGISTERS_4_18_port, ZN => n14718);
   U12923 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_18_port, B1 => 
                           n15119, B2 => REGISTERS_7_18_port, ZN => n14717);
   U12924 : AND4_X1 port map( A1 => n14720, A2 => n14719, A3 => n14718, A4 => 
                           n14717, ZN => n14737);
   U12925 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_18_port, B1 => 
                           n15142, B2 => REGISTERS_14_18_port, ZN => n14724);
   U12926 : AOI22_X1 port map( A1 => n15145, A2 => REGISTERS_8_18_port, B1 => 
                           n15144, B2 => REGISTERS_9_18_port, ZN => n14723);
   U12927 : AOI22_X1 port map( A1 => n15033, A2 => REGISTERS_26_18_port, B1 => 
                           n15130, B2 => REGISTERS_16_18_port, ZN => n14722);
   U12928 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_18_port, B1 => 
                           n15128, B2 => REGISTERS_22_18_port, ZN => n14721);
   U12929 : NAND4_X1 port map( A1 => n14724, A2 => n14723, A3 => n14722, A4 => 
                           n14721, ZN => n14735);
   U12930 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_18_port, B1 => 
                           n15154, B2 => REGISTERS_21_18_port, ZN => n14728);
   U12931 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_18_port, B1 => 
                           n15156, B2 => REGISTERS_23_18_port, ZN => n14727);
   U12932 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_18_port, B1 => 
                           n15133, B2 => REGISTERS_30_18_port, ZN => n14726);
   U12933 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_18_port, B1 => 
                           n15151, B2 => REGISTERS_28_18_port, ZN => n14725);
   U12934 : NAND4_X1 port map( A1 => n14728, A2 => n14727, A3 => n14726, A4 => 
                           n14725, ZN => n14734);
   U12935 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_18_port, B1 => 
                           n15127, B2 => REGISTERS_24_18_port, ZN => n14732);
   U12936 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_18_port, B1 => 
                           n15155, B2 => REGISTERS_18_18_port, ZN => n14731);
   U12937 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_18_port, B1 => 
                           n15150, B2 => REGISTERS_10_18_port, ZN => n14730);
   U12938 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_18_port, B1 => 
                           n15126, B2 => REGISTERS_29_18_port, ZN => n14729);
   U12939 : NAND4_X1 port map( A1 => n14732, A2 => n14731, A3 => n14730, A4 => 
                           n14729, ZN => n14733);
   U12940 : NOR3_X1 port map( A1 => n14735, A2 => n14734, A3 => n14733, ZN => 
                           n14736);
   U12941 : OAI222_X1 port map( A1 => n14910, A2 => n8460, B1 => n14505, B2 => 
                           n14737, C1 => n14354, C2 => n14736, ZN => n8551);
   U12942 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_17_port, B1 => 
                           n15119, B2 => REGISTERS_7_17_port, ZN => n14741);
   U12943 : AOI22_X1 port map( A1 => n14483, A2 => REGISTERS_4_17_port, B1 => 
                           n15116, B2 => REGISTERS_0_17_port, ZN => n14740);
   U12944 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_17_port, B1 => 
                           n14781, B2 => REGISTERS_6_17_port, ZN => n14739);
   U12945 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_17_port, B1 => 
                           n15088, B2 => REGISTERS_5_17_port, ZN => n14738);
   U12946 : AND4_X1 port map( A1 => n14741, A2 => n14740, A3 => n14739, A4 => 
                           n14738, ZN => n14758);
   U12947 : AOI22_X1 port map( A1 => n15033, A2 => REGISTERS_26_17_port, B1 => 
                           n15154, B2 => REGISTERS_21_17_port, ZN => n14745);
   U12948 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_17_port, B1 => 
                           n15152, B2 => REGISTERS_31_17_port, ZN => n14744);
   U12949 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_17_port, B1 => 
                           n15126, B2 => REGISTERS_29_17_port, ZN => n14743);
   U12950 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_17_port, B1 => 
                           n15138, B2 => REGISTERS_11_17_port, ZN => n14742);
   U12951 : NAND4_X1 port map( A1 => n14745, A2 => n14744, A3 => n14743, A4 => 
                           n14742, ZN => n14756);
   U12952 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_17_port, B1 => 
                           n15128, B2 => REGISTERS_22_17_port, ZN => n14749);
   U12953 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_17_port, B1 => 
                           n15096, B2 => REGISTERS_28_17_port, ZN => n14748);
   U12954 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_17_port, B1 => 
                           n15139, B2 => REGISTERS_19_17_port, ZN => n14747);
   U12955 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_17_port, B1 => 
                           n15144, B2 => REGISTERS_9_17_port, ZN => n14746);
   U12956 : NAND4_X1 port map( A1 => n14749, A2 => n14748, A3 => n14747, A4 => 
                           n14746, ZN => n14755);
   U12957 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_17_port, B1 => 
                           n15130, B2 => REGISTERS_16_17_port, ZN => n14753);
   U12958 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_17_port, B1 => 
                           n15132, B2 => REGISTERS_15_17_port, ZN => n14752);
   U12959 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_17_port, B1 => 
                           n15145, B2 => REGISTERS_8_17_port, ZN => n14751);
   U12960 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_17_port, B1 => 
                           n15142, B2 => REGISTERS_14_17_port, ZN => n14750);
   U12961 : NAND4_X1 port map( A1 => n14753, A2 => n14752, A3 => n14751, A4 => 
                           n14750, ZN => n14754);
   U12962 : NOR3_X1 port map( A1 => n14756, A2 => n14755, A3 => n14754, ZN => 
                           n14757);
   U12963 : OAI222_X1 port map( A1 => n16071, A2 => n8459, B1 => n15115, B2 => 
                           n14758, C1 => n15166, C2 => n14757, ZN => n8552);
   U12964 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_16_port, B1 => 
                           n15116, B2 => REGISTERS_0_16_port, ZN => n14763);
   U12965 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_16_port, B1 => 
                           n15091, B2 => REGISTERS_7_16_port, ZN => n14762);
   U12966 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_16_port, B1 => 
                           n14781, B2 => REGISTERS_6_16_port, ZN => n14761);
   U12967 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_16_port, B1 => 
                           n14483, B2 => REGISTERS_4_16_port, ZN => n14760);
   U12968 : AND4_X1 port map( A1 => n14763, A2 => n14762, A3 => n14761, A4 => 
                           n14760, ZN => n14780);
   U12969 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_16_port, B1 => 
                           n15143, B2 => REGISTERS_27_16_port, ZN => n14767);
   U12970 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_16_port, B1 => 
                           n15128, B2 => REGISTERS_22_16_port, ZN => n14766);
   U12971 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_16_port, B1 => 
                           n15154, B2 => REGISTERS_21_16_port, ZN => n14765);
   U12972 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_16_port, B1 => 
                           n15144, B2 => REGISTERS_9_16_port, ZN => n14764);
   U12973 : NAND4_X1 port map( A1 => n14767, A2 => n14766, A3 => n14765, A4 => 
                           n14764, ZN => n14778);
   U12974 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_16_port, B1 => 
                           n15126, B2 => REGISTERS_29_16_port, ZN => n14771);
   U12975 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_16_port, B1 => 
                           n14944, B2 => REGISTERS_25_16_port, ZN => n14770);
   U12976 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_16_port, B1 => 
                           n15130, B2 => REGISTERS_16_16_port, ZN => n14769);
   U12977 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_16_port, B1 => 
                           n15150, B2 => REGISTERS_10_16_port, ZN => n14768);
   U12978 : NAND4_X1 port map( A1 => n14771, A2 => n14770, A3 => n14769, A4 => 
                           n14768, ZN => n14777);
   U12979 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_16_port, B1 => 
                           n15153, B2 => REGISTERS_20_16_port, ZN => n14775);
   U12980 : AOI22_X1 port map( A1 => n15142, A2 => REGISTERS_14_16_port, B1 => 
                           n15145, B2 => REGISTERS_8_16_port, ZN => n14774);
   U12981 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_16_port, B1 => 
                           n14837, B2 => REGISTERS_28_16_port, ZN => n14773);
   U12982 : AOI22_X1 port map( A1 => n15033, A2 => REGISTERS_26_16_port, B1 => 
                           n15129, B2 => REGISTERS_17_16_port, ZN => n14772);
   U12983 : NAND4_X1 port map( A1 => n14775, A2 => n14774, A3 => n14773, A4 => 
                           n14772, ZN => n14776);
   U12984 : NOR3_X1 port map( A1 => n14778, A2 => n14777, A3 => n14776, ZN => 
                           n14779);
   U12985 : OAI222_X1 port map( A1 => n16071, A2 => n8458, B1 => n14505, B2 => 
                           n14780, C1 => n14354, C2 => n14779, ZN => n8553);
   U12986 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_15_port, B1 => 
                           n14781, B2 => REGISTERS_6_15_port, ZN => n14785);
   U12987 : AOI22_X1 port map( A1 => n15117, A2 => REGISTERS_4_15_port, B1 => 
                           n15089, B2 => REGISTERS_0_15_port, ZN => n14784);
   U12988 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_15_port, B1 => 
                           n15091, B2 => REGISTERS_7_15_port, ZN => n14783);
   U12989 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_15_port, B1 => 
                           n15088, B2 => REGISTERS_5_15_port, ZN => n14782);
   U12990 : AND4_X1 port map( A1 => n14785, A2 => n14784, A3 => n14783, A4 => 
                           n14782, ZN => n14802);
   U12991 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_15_port, B1 => 
                           n15133, B2 => REGISTERS_30_15_port, ZN => n14789);
   U12992 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_15_port, B1 => 
                           n15152, B2 => REGISTERS_31_15_port, ZN => n14788);
   U12993 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_15_port, B1 => 
                           n15150, B2 => REGISTERS_10_15_port, ZN => n14787);
   U12994 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_15_port, B1 => 
                           n15156, B2 => REGISTERS_23_15_port, ZN => n14786);
   U12995 : NAND4_X1 port map( A1 => n14789, A2 => n14788, A3 => n14787, A4 => 
                           n14786, ZN => n14800);
   U12996 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_15_port, B1 => 
                           n15154, B2 => REGISTERS_21_15_port, ZN => n14793);
   U12997 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_15_port, B1 => 
                           n15138, B2 => REGISTERS_11_15_port, ZN => n14792);
   U12998 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_15_port, B1 => 
                           n15130, B2 => REGISTERS_16_15_port, ZN => n14791);
   U12999 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_15_port, B1 => 
                           n15127, B2 => REGISTERS_24_15_port, ZN => n14790);
   U13000 : NAND4_X1 port map( A1 => n14793, A2 => n14792, A3 => n14791, A4 => 
                           n14790, ZN => n14799);
   U13001 : AOI22_X1 port map( A1 => n15096, A2 => REGISTERS_28_15_port, B1 => 
                           n15144, B2 => REGISTERS_9_15_port, ZN => n14797);
   U13002 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_15_port, B1 => 
                           n15145, B2 => REGISTERS_8_15_port, ZN => n14796);
   U13003 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_15_port, B1 => 
                           n15142, B2 => REGISTERS_14_15_port, ZN => n14795);
   U13004 : AOI22_X1 port map( A1 => n15126, A2 => REGISTERS_29_15_port, B1 => 
                           n15128, B2 => REGISTERS_22_15_port, ZN => n14794);
   U13005 : NAND4_X1 port map( A1 => n14797, A2 => n14796, A3 => n14795, A4 => 
                           n14794, ZN => n14798);
   U13006 : NOR3_X1 port map( A1 => n14800, A2 => n14799, A3 => n14798, ZN => 
                           n14801);
   U13007 : OAI222_X1 port map( A1 => n16026, A2 => n8457, B1 => n15115, B2 => 
                           n14802, C1 => n15166, C2 => n14801, ZN => n8554);
   U13008 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_14_port, B1 => 
                           n15117, B2 => REGISTERS_4_14_port, ZN => n14806);
   U13009 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_14_port, B1 => 
                           n15121, B2 => REGISTERS_3_14_port, ZN => n14805);
   U13010 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_14_port, B1 => 
                           n15119, B2 => REGISTERS_7_14_port, ZN => n14804);
   U13011 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_14_port, B1 => 
                           n15089, B2 => REGISTERS_0_14_port, ZN => n14803);
   U13012 : AND4_X1 port map( A1 => n14806, A2 => n14805, A3 => n14804, A4 => 
                           n14803, ZN => n14823);
   U13013 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_14_port, B1 => 
                           n15157, B2 => REGISTERS_13_14_port, ZN => n14810);
   U13014 : AOI22_X1 port map( A1 => n15142, A2 => REGISTERS_14_14_port, B1 => 
                           n15154, B2 => REGISTERS_21_14_port, ZN => n14809);
   U13015 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_14_port, B1 => 
                           n15150, B2 => REGISTERS_10_14_port, ZN => n14808);
   U13016 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_14_port, B1 => 
                           n15132, B2 => REGISTERS_15_14_port, ZN => n14807);
   U13017 : NAND4_X1 port map( A1 => n14810, A2 => n14809, A3 => n14808, A4 => 
                           n14807, ZN => n14821);
   U13018 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_14_port, B1 => 
                           n15138, B2 => REGISTERS_11_14_port, ZN => n14814);
   U13019 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_14_port, B1 => 
                           n15152, B2 => REGISTERS_31_14_port, ZN => n14813);
   U13020 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_14_port, B1 => 
                           n15151, B2 => REGISTERS_28_14_port, ZN => n14812);
   U13021 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_14_port, B1 => 
                           n15143, B2 => REGISTERS_27_14_port, ZN => n14811);
   U13022 : NAND4_X1 port map( A1 => n14814, A2 => n14813, A3 => n14812, A4 => 
                           n14811, ZN => n14820);
   U13023 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_14_port, B1 => 
                           n15144, B2 => REGISTERS_9_14_port, ZN => n14818);
   U13024 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_14_port, B1 => 
                           n15130, B2 => REGISTERS_16_14_port, ZN => n14817);
   U13025 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_14_port, B1 => 
                           n15126, B2 => REGISTERS_29_14_port, ZN => n14816);
   U13026 : AOI22_X1 port map( A1 => n15145, A2 => REGISTERS_8_14_port, B1 => 
                           n15128, B2 => REGISTERS_22_14_port, ZN => n14815);
   U13027 : NAND4_X1 port map( A1 => n14818, A2 => n14817, A3 => n14816, A4 => 
                           n14815, ZN => n14819);
   U13028 : NOR3_X1 port map( A1 => n14821, A2 => n14820, A3 => n14819, ZN => 
                           n14822);
   U13029 : OAI222_X1 port map( A1 => n14910, A2 => n8456, B1 => n15115, B2 => 
                           n14823, C1 => n14354, C2 => n14822, ZN => n8555);
   U13030 : AOI22_X1 port map( A1 => n15091, A2 => REGISTERS_7_13_port, B1 => 
                           n15116, B2 => REGISTERS_0_13_port, ZN => n14827);
   U13031 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_13_port, B1 => 
                           n14483, B2 => REGISTERS_4_13_port, ZN => n14826);
   U13032 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_13_port, B1 => 
                           n15088, B2 => REGISTERS_5_13_port, ZN => n14825);
   U13033 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_13_port, B1 => 
                           n15121, B2 => REGISTERS_3_13_port, ZN => n14824);
   U13034 : AND4_X1 port map( A1 => n14827, A2 => n14826, A3 => n14825, A4 => 
                           n14824, ZN => n14846);
   U13035 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_13_port, B1 => 
                           n15126, B2 => REGISTERS_29_13_port, ZN => n14831);
   U13036 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_13_port, B1 => 
                           n15154, B2 => REGISTERS_21_13_port, ZN => n14830);
   U13037 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_13_port, B1 => 
                           n15032, B2 => REGISTERS_30_13_port, ZN => n14829);
   U13038 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_13_port, B1 => 
                           n15140, B2 => REGISTERS_12_13_port, ZN => n14828);
   U13039 : NAND4_X1 port map( A1 => n14831, A2 => n14830, A3 => n14829, A4 => 
                           n14828, ZN => n14844);
   U13040 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_13_port, B1 => 
                           n15142, B2 => REGISTERS_14_13_port, ZN => n14836);
   U13041 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_13_port, B1 => 
                           n15145, B2 => REGISTERS_8_13_port, ZN => n14835);
   U13042 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_13_port, B1 => 
                           n15144, B2 => REGISTERS_9_13_port, ZN => n14834);
   U13043 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_13_port, B1 => 
                           n15130, B2 => REGISTERS_16_13_port, ZN => n14833);
   U13044 : NAND4_X1 port map( A1 => n14836, A2 => n14835, A3 => n14834, A4 => 
                           n14833, ZN => n14843);
   U13045 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_13_port, B1 => 
                           n15143, B2 => REGISTERS_27_13_port, ZN => n14841);
   U13046 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_13_port, B1 => 
                           n15127, B2 => REGISTERS_24_13_port, ZN => n14840);
   U13047 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_13_port, B1 => 
                           n15128, B2 => REGISTERS_22_13_port, ZN => n14839);
   U13048 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_13_port, B1 => 
                           n14837, B2 => REGISTERS_28_13_port, ZN => n14838);
   U13049 : NAND4_X1 port map( A1 => n14841, A2 => n14840, A3 => n14839, A4 => 
                           n14838, ZN => n14842);
   U13050 : NOR3_X1 port map( A1 => n14844, A2 => n14843, A3 => n14842, ZN => 
                           n14845);
   U13051 : OAI222_X1 port map( A1 => n16071, A2 => n8455, B1 => n15115, B2 => 
                           n14846, C1 => n15166, C2 => n14845, ZN => n8556);
   U13052 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_12_port, B1 => 
                           n15116, B2 => REGISTERS_0_12_port, ZN => n14850);
   U13053 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_12_port, B1 => 
                           n14483, B2 => REGISTERS_4_12_port, ZN => n14849);
   U13054 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_12_port, B1 => 
                           n15120, B2 => REGISTERS_1_12_port, ZN => n14848);
   U13055 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_12_port, B1 => 
                           n15091, B2 => REGISTERS_7_12_port, ZN => n14847);
   U13056 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_12_port, B1 => 
                           n15156, B2 => REGISTERS_23_12_port, ZN => n14854);
   U13057 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_12_port, B1 => 
                           n15150, B2 => REGISTERS_10_12_port, ZN => n14853);
   U13058 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_12_port, B1 => 
                           n15154, B2 => REGISTERS_21_12_port, ZN => n14852);
   U13059 : AOI22_X1 port map( A1 => n15096, A2 => REGISTERS_28_12_port, B1 => 
                           n15128, B2 => REGISTERS_22_12_port, ZN => n14851);
   U13060 : NAND4_X1 port map( A1 => n14854, A2 => n14853, A3 => n14852, A4 => 
                           n14851, ZN => n14865);
   U13061 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_12_port, B1 => 
                           n15155, B2 => REGISTERS_18_12_port, ZN => n14858);
   U13062 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_12_port, B1 => 
                           n14979, B2 => REGISTERS_19_12_port, ZN => n14857);
   U13063 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_12_port, B1 => 
                           n15130, B2 => REGISTERS_16_12_port, ZN => n14856);
   U13064 : AOI22_X1 port map( A1 => n15144, A2 => REGISTERS_9_12_port, B1 => 
                           n15126, B2 => REGISTERS_29_12_port, ZN => n14855);
   U13065 : NAND4_X1 port map( A1 => n14858, A2 => n14857, A3 => n14856, A4 => 
                           n14855, ZN => n14864);
   U13066 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_12_port, B1 => 
                           n15127, B2 => REGISTERS_24_12_port, ZN => n14862);
   U13067 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_12_port, B1 => 
                           n15145, B2 => REGISTERS_8_12_port, ZN => n14861);
   U13068 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_12_port, B1 => 
                           n15142, B2 => REGISTERS_14_12_port, ZN => n14860);
   U13069 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_12_port, B1 => 
                           n15132, B2 => REGISTERS_15_12_port, ZN => n14859);
   U13070 : NAND4_X1 port map( A1 => n14862, A2 => n14861, A3 => n14860, A4 => 
                           n14859, ZN => n14863);
   U13071 : NOR3_X1 port map( A1 => n14865, A2 => n14864, A3 => n14863, ZN => 
                           n14866);
   U13072 : OAI222_X1 port map( A1 => n14910, A2 => n8454, B1 => n14505, B2 => 
                           n14867, C1 => n14354, C2 => n14866, ZN => n8557);
   U13073 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_11_port, B1 => 
                           n14483, B2 => REGISTERS_4_11_port, ZN => n14871);
   U13074 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_11_port, B1 => 
                           n15089, B2 => REGISTERS_0_11_port, ZN => n14870);
   U13075 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_11_port, B1 => 
                           n15088, B2 => REGISTERS_5_11_port, ZN => n14869);
   U13076 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_11_port, B1 => 
                           n15119, B2 => REGISTERS_7_11_port, ZN => n14868);
   U13077 : AND4_X1 port map( A1 => n14871, A2 => n14870, A3 => n14869, A4 => 
                           n14868, ZN => n14888);
   U13078 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_11_port, B1 => 
                           n15154, B2 => REGISTERS_21_11_port, ZN => n14875);
   U13079 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_11_port, B1 => 
                           n15145, B2 => REGISTERS_8_11_port, ZN => n14874);
   U13080 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_11_port, B1 => 
                           n15096, B2 => REGISTERS_28_11_port, ZN => n14873);
   U13081 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_11_port, B1 => 
                           n15144, B2 => REGISTERS_9_11_port, ZN => n14872);
   U13082 : NAND4_X1 port map( A1 => n14875, A2 => n14874, A3 => n14873, A4 => 
                           n14872, ZN => n14886);
   U13083 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_11_port, B1 => 
                           n15132, B2 => REGISTERS_15_11_port, ZN => n14879);
   U13084 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_11_port, B1 => 
                           n15126, B2 => REGISTERS_29_11_port, ZN => n14878);
   U13085 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_11_port, B1 => 
                           n15141, B2 => REGISTERS_25_11_port, ZN => n14877);
   U13086 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_11_port, B1 => 
                           n15127, B2 => REGISTERS_24_11_port, ZN => n14876);
   U13087 : NAND4_X1 port map( A1 => n14879, A2 => n14878, A3 => n14877, A4 => 
                           n14876, ZN => n14885);
   U13088 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_11_port, B1 => 
                           n15128, B2 => REGISTERS_22_11_port, ZN => n14883);
   U13089 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_11_port, B1 => 
                           n15156, B2 => REGISTERS_23_11_port, ZN => n14882);
   U13090 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_11_port, B1 => 
                           n15142, B2 => REGISTERS_14_11_port, ZN => n14881);
   U13091 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_11_port, B1 => 
                           n15130, B2 => REGISTERS_16_11_port, ZN => n14880);
   U13092 : NAND4_X1 port map( A1 => n14883, A2 => n14882, A3 => n14881, A4 => 
                           n14880, ZN => n14884);
   U13093 : NOR3_X1 port map( A1 => n14886, A2 => n14885, A3 => n14884, ZN => 
                           n14887);
   U13094 : OAI222_X1 port map( A1 => n16026, A2 => n8453, B1 => n15115, B2 => 
                           n14888, C1 => n14354, C2 => n14887, ZN => n8558);
   U13095 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_10_port, B1 => 
                           n15117, B2 => REGISTERS_4_10_port, ZN => n14892);
   U13096 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_10_port, B1 => 
                           n15043, B2 => REGISTERS_6_10_port, ZN => n14891);
   U13097 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_10_port, B1 => 
                           n15120, B2 => REGISTERS_1_10_port, ZN => n14890);
   U13098 : AOI22_X1 port map( A1 => n15091, A2 => REGISTERS_7_10_port, B1 => 
                           n15116, B2 => REGISTERS_0_10_port, ZN => n14889);
   U13099 : AND4_X1 port map( A1 => n14892, A2 => n14891, A3 => n14890, A4 => 
                           n14889, ZN => n14909);
   U13100 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_10_port, B1 => 
                           n15096, B2 => REGISTERS_28_10_port, ZN => n14896);
   U13101 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_10_port, B1 => 
                           n15145, B2 => REGISTERS_8_10_port, ZN => n14895);
   U13102 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_10_port, B1 => 
                           n15156, B2 => REGISTERS_23_10_port, ZN => n14894);
   U13103 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_10_port, B1 => 
                           n15153, B2 => REGISTERS_20_10_port, ZN => n14893);
   U13104 : NAND4_X1 port map( A1 => n14896, A2 => n14895, A3 => n14894, A4 => 
                           n14893, ZN => n14907);
   U13105 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_10_port, B1 => 
                           n14944, B2 => REGISTERS_25_10_port, ZN => n14900);
   U13106 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_10_port, B1 => 
                           n15144, B2 => REGISTERS_9_10_port, ZN => n14899);
   U13107 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_10_port, B1 => 
                           n15032, B2 => REGISTERS_30_10_port, ZN => n14898);
   U13108 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_10_port, B1 => 
                           n15132, B2 => REGISTERS_15_10_port, ZN => n14897);
   U13109 : NAND4_X1 port map( A1 => n14900, A2 => n14899, A3 => n14898, A4 => 
                           n14897, ZN => n14906);
   U13110 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_10_port, B1 => 
                           n15154, B2 => REGISTERS_21_10_port, ZN => n14904);
   U13111 : AOI22_X1 port map( A1 => n15126, A2 => REGISTERS_29_10_port, B1 => 
                           n15128, B2 => REGISTERS_22_10_port, ZN => n14903);
   U13112 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_10_port, B1 => 
                           n15150, B2 => REGISTERS_10_10_port, ZN => n14902);
   U13113 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_10_port, B1 => 
                           n15142, B2 => REGISTERS_14_10_port, ZN => n14901);
   U13114 : NAND4_X1 port map( A1 => n14904, A2 => n14903, A3 => n14902, A4 => 
                           n14901, ZN => n14905);
   U13115 : NOR3_X1 port map( A1 => n14907, A2 => n14906, A3 => n14905, ZN => 
                           n14908);
   U13116 : OAI222_X1 port map( A1 => n14910, A2 => n8452, B1 => n15115, B2 => 
                           n14909, C1 => n15166, C2 => n14908, ZN => n8559);
   U13117 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_9_port, B1 => 
                           n15091, B2 => REGISTERS_7_9_port, ZN => n14914);
   U13118 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_9_port, B1 => 
                           n15117, B2 => REGISTERS_4_9_port, ZN => n14913);
   U13119 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_9_port, B1 => 
                           n15090, B2 => REGISTERS_3_9_port, ZN => n14912);
   U13120 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_9_port, B1 => 
                           n15089, B2 => REGISTERS_0_9_port, ZN => n14911);
   U13121 : AND4_X1 port map( A1 => n14914, A2 => n14913, A3 => n14912, A4 => 
                           n14911, ZN => n14931);
   U13122 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_9_port, B1 => 
                           n15154, B2 => REGISTERS_21_9_port, ZN => n14918);
   U13123 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_9_port, B1 => 
                           n15144, B2 => REGISTERS_9_9_port, ZN => n14917);
   U13124 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_9_port, B1 => 
                           n15140, B2 => REGISTERS_12_9_port, ZN => n14916);
   U13125 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_9_port, B1 => 
                           n15142, B2 => REGISTERS_14_9_port, ZN => n14915);
   U13126 : NAND4_X1 port map( A1 => n14918, A2 => n14917, A3 => n14916, A4 => 
                           n14915, ZN => n14929);
   U13127 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_9_port, B1 => 
                           n15127, B2 => REGISTERS_24_9_port, ZN => n14922);
   U13128 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_9_port, B1 => 
                           n15096, B2 => REGISTERS_28_9_port, ZN => n14921);
   U13129 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_9_port, B1 => 
                           n15150, B2 => REGISTERS_10_9_port, ZN => n14920);
   U13130 : AOI22_X1 port map( A1 => n15145, A2 => REGISTERS_8_9_port, B1 => 
                           n15128, B2 => REGISTERS_22_9_port, ZN => n14919);
   U13131 : NAND4_X1 port map( A1 => n14922, A2 => n14921, A3 => n14920, A4 => 
                           n14919, ZN => n14928);
   U13132 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_9_port, B1 => 
                           n15156, B2 => REGISTERS_23_9_port, ZN => n14926);
   U13133 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_9_port, B1 => 
                           n15153, B2 => REGISTERS_20_9_port, ZN => n14925);
   U13134 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_9_port, B1 => 
                           n15126, B2 => REGISTERS_29_9_port, ZN => n14924);
   U13135 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_9_port, B1 => 
                           n15132, B2 => REGISTERS_15_9_port, ZN => n14923);
   U13136 : NAND4_X1 port map( A1 => n14926, A2 => n14925, A3 => n14924, A4 => 
                           n14923, ZN => n14927);
   U13137 : NOR3_X1 port map( A1 => n14929, A2 => n14928, A3 => n14927, ZN => 
                           n14930);
   U13138 : OAI222_X1 port map( A1 => n16071, A2 => n8451, B1 => n15115, B2 => 
                           n14931, C1 => n14354, C2 => n14930, ZN => n8560);
   U13139 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_8_port, B1 => 
                           n14483, B2 => REGISTERS_4_8_port, ZN => n14935);
   U13140 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_8_port, B1 => 
                           n15116, B2 => REGISTERS_0_8_port, ZN => n14934);
   U13141 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_8_port, B1 => 
                           n15119, B2 => REGISTERS_7_8_port, ZN => n14933);
   U13142 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_8_port, B1 => 
                           n15043, B2 => REGISTERS_6_8_port, ZN => n14932);
   U13143 : AND4_X1 port map( A1 => n14935, A2 => n14934, A3 => n14933, A4 => 
                           n14932, ZN => n14953);
   U13144 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_8_port, B1 => 
                           n15143, B2 => REGISTERS_27_8_port, ZN => n14939);
   U13145 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_8_port, B1 => 
                           n15153, B2 => REGISTERS_20_8_port, ZN => n14938);
   U13146 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_8_port, B1 => 
                           n15129, B2 => REGISTERS_17_8_port, ZN => n14937);
   U13147 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_8_port, B1 => 
                           n15145, B2 => REGISTERS_8_8_port, ZN => n14936);
   U13148 : NAND4_X1 port map( A1 => n14939, A2 => n14938, A3 => n14937, A4 => 
                           n14936, ZN => n14951);
   U13149 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_8_port, B1 => 
                           n15128, B2 => REGISTERS_22_8_port, ZN => n14943);
   U13150 : AOI22_X1 port map( A1 => n15126, A2 => REGISTERS_29_8_port, B1 => 
                           n15154, B2 => REGISTERS_21_8_port, ZN => n14942);
   U13151 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_8_port, B1 => 
                           n15156, B2 => REGISTERS_23_8_port, ZN => n14941);
   U13152 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_8_port, B1 => 
                           n15142, B2 => REGISTERS_14_8_port, ZN => n14940);
   U13153 : NAND4_X1 port map( A1 => n14943, A2 => n14942, A3 => n14941, A4 => 
                           n14940, ZN => n14950);
   U13154 : AOI22_X1 port map( A1 => n14944, A2 => REGISTERS_25_8_port, B1 => 
                           n15151, B2 => REGISTERS_28_8_port, ZN => n14948);
   U13155 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_8_port, B1 => 
                           n15150, B2 => REGISTERS_10_8_port, ZN => n14947);
   U13156 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_8_port, B1 => 
                           n15144, B2 => REGISTERS_9_8_port, ZN => n14946);
   U13157 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_8_port, B1 => 
                           n15152, B2 => REGISTERS_31_8_port, ZN => n14945);
   U13158 : NAND4_X1 port map( A1 => n14948, A2 => n14947, A3 => n14946, A4 => 
                           n14945, ZN => n14949);
   U13159 : NOR3_X1 port map( A1 => n14951, A2 => n14950, A3 => n14949, ZN => 
                           n14952);
   U13160 : OAI222_X1 port map( A1 => n16071, A2 => n8450, B1 => n14505, B2 => 
                           n14953, C1 => n15166, C2 => n14952, ZN => n8561);
   U13161 : AOI22_X1 port map( A1 => n15117, A2 => REGISTERS_4_7_port, B1 => 
                           n15091, B2 => REGISTERS_7_7_port, ZN => n14957);
   U13162 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_7_port, B1 => 
                           n15089, B2 => REGISTERS_0_7_port, ZN => n14956);
   U13163 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_7_port, B1 => 
                           n15088, B2 => REGISTERS_5_7_port, ZN => n14955);
   U13164 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_7_port, B1 => 
                           n15090, B2 => REGISTERS_3_7_port, ZN => n14954);
   U13165 : AND4_X1 port map( A1 => n14957, A2 => n14956, A3 => n14955, A4 => 
                           n14954, ZN => n14974);
   U13166 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_7_port, B1 => 
                           n15140, B2 => REGISTERS_12_7_port, ZN => n14961);
   U13167 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_7_port, B1 => 
                           n15132, B2 => REGISTERS_15_7_port, ZN => n14960);
   U13168 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_7_port, B1 => 
                           n15154, B2 => REGISTERS_21_7_port, ZN => n14959);
   U13169 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_7_port, B1 => 
                           n15130, B2 => REGISTERS_16_7_port, ZN => n14958);
   U13170 : NAND4_X1 port map( A1 => n14961, A2 => n14960, A3 => n14959, A4 => 
                           n14958, ZN => n14972);
   U13171 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_7_port, B1 => 
                           n15126, B2 => REGISTERS_29_7_port, ZN => n14965);
   U13172 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_7_port, B1 => 
                           n15155, B2 => REGISTERS_18_7_port, ZN => n14964);
   U13173 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_7_port, B1 => 
                           n15096, B2 => REGISTERS_28_7_port, ZN => n14963);
   U13174 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_7_port, B1 => 
                           n15142, B2 => REGISTERS_14_7_port, ZN => n14962);
   U13175 : NAND4_X1 port map( A1 => n14965, A2 => n14964, A3 => n14963, A4 => 
                           n14962, ZN => n14971);
   U13176 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_7_port, B1 => 
                           n15144, B2 => REGISTERS_9_7_port, ZN => n14969);
   U13177 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_7_port, B1 => 
                           n15128, B2 => REGISTERS_22_7_port, ZN => n14968);
   U13178 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_7_port, B1 => 
                           n15145, B2 => REGISTERS_8_7_port, ZN => n14967);
   U13179 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_7_port, B1 => 
                           n15150, B2 => REGISTERS_10_7_port, ZN => n14966);
   U13180 : NAND4_X1 port map( A1 => n14969, A2 => n14968, A3 => n14967, A4 => 
                           n14966, ZN => n14970);
   U13181 : NOR3_X1 port map( A1 => n14972, A2 => n14971, A3 => n14970, ZN => 
                           n14973);
   U13182 : OAI222_X1 port map( A1 => n16026, A2 => n8449, B1 => n15115, B2 => 
                           n14974, C1 => n14354, C2 => n14973, ZN => n8562);
   U13183 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_6_port, B1 => 
                           n15043, B2 => REGISTERS_6_6_port, ZN => n14978);
   U13184 : AOI22_X1 port map( A1 => n14483, A2 => REGISTERS_4_6_port, B1 => 
                           n15089, B2 => REGISTERS_0_6_port, ZN => n14977);
   U13185 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_6_port, B1 => 
                           n15119, B2 => REGISTERS_7_6_port, ZN => n14976);
   U13186 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_6_port, B1 => 
                           n15090, B2 => REGISTERS_3_6_port, ZN => n14975);
   U13187 : AND4_X1 port map( A1 => n14978, A2 => n14977, A3 => n14976, A4 => 
                           n14975, ZN => n14996);
   U13188 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_6_port, B1 => 
                           n15126, B2 => REGISTERS_29_6_port, ZN => n14983);
   U13189 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_6_port, B1 => 
                           n15154, B2 => REGISTERS_21_6_port, ZN => n14982);
   U13190 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_6_port, B1 => 
                           n14979, B2 => REGISTERS_19_6_port, ZN => n14981);
   U13191 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_6_port, B1 => 
                           n15152, B2 => REGISTERS_31_6_port, ZN => n14980);
   U13192 : NAND4_X1 port map( A1 => n14983, A2 => n14982, A3 => n14981, A4 => 
                           n14980, ZN => n14994);
   U13193 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_6_port, B1 => 
                           n15128, B2 => REGISTERS_22_6_port, ZN => n14987);
   U13194 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_6_port, B1 => 
                           n15130, B2 => REGISTERS_16_6_port, ZN => n14986);
   U13195 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_6_port, B1 => 
                           n15138, B2 => REGISTERS_11_6_port, ZN => n14985);
   U13196 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_6_port, B1 => 
                           n15144, B2 => REGISTERS_9_6_port, ZN => n14984);
   U13197 : NAND4_X1 port map( A1 => n14987, A2 => n14986, A3 => n14985, A4 => 
                           n14984, ZN => n14993);
   U13198 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_6_port, B1 => 
                           n15145, B2 => REGISTERS_8_6_port, ZN => n14991);
   U13199 : AOI22_X1 port map( A1 => n15140, A2 => REGISTERS_12_6_port, B1 => 
                           n15151, B2 => REGISTERS_28_6_port, ZN => n14990);
   U13200 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_6_port, B1 => 
                           n15142, B2 => REGISTERS_14_6_port, ZN => n14989);
   U13201 : AOI22_X1 port map( A1 => n15074, A2 => REGISTERS_30_6_port, B1 => 
                           n15150, B2 => REGISTERS_10_6_port, ZN => n14988);
   U13202 : NAND4_X1 port map( A1 => n14991, A2 => n14990, A3 => n14989, A4 => 
                           n14988, ZN => n14992);
   U13203 : NOR3_X1 port map( A1 => n14994, A2 => n14993, A3 => n14992, ZN => 
                           n14995);
   U13204 : OAI222_X1 port map( A1 => n16071, A2 => n8448, B1 => n15115, B2 => 
                           n14996, C1 => n15166, C2 => n14995, ZN => n8563);
   U13205 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_5_port, B1 => 
                           n15116, B2 => REGISTERS_0_5_port, ZN => n15000);
   U13206 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_5_port, B1 => 
                           n15091, B2 => REGISTERS_7_5_port, ZN => n14999);
   U13207 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_5_port, B1 => 
                           n15120, B2 => REGISTERS_1_5_port, ZN => n14998);
   U13208 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_5_port, B1 => 
                           n15117, B2 => REGISTERS_4_5_port, ZN => n14997);
   U13209 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_5_port, B1 => 
                           n15144, B2 => REGISTERS_9_5_port, ZN => n15004);
   U13210 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_5_port, B1 => 
                           n15128, B2 => REGISTERS_22_5_port, ZN => n15003);
   U13211 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_5_port, B1 => 
                           n15142, B2 => REGISTERS_14_5_port, ZN => n15002);
   U13212 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_5_port, B1 => 
                           n15130, B2 => REGISTERS_16_5_port, ZN => n15001);
   U13213 : NAND4_X1 port map( A1 => n15004, A2 => n15003, A3 => n15002, A4 => 
                           n15001, ZN => n15016);
   U13214 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_5_port, B1 => 
                           n15156, B2 => REGISTERS_23_5_port, ZN => n15009);
   U13215 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_5_port, B1 => 
                           n15140, B2 => REGISTERS_12_5_port, ZN => n15008);
   U13216 : AOI22_X1 port map( A1 => n15005, A2 => REGISTERS_26_5_port, B1 => 
                           n15129, B2 => REGISTERS_17_5_port, ZN => n15007);
   U13217 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_5_port, B1 => 
                           n15126, B2 => REGISTERS_29_5_port, ZN => n15006);
   U13218 : NAND4_X1 port map( A1 => n15009, A2 => n15008, A3 => n15007, A4 => 
                           n15006, ZN => n15015);
   U13219 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_5_port, B1 => 
                           n15096, B2 => REGISTERS_28_5_port, ZN => n15013);
   U13220 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_5_port, B1 => 
                           n15132, B2 => REGISTERS_15_5_port, ZN => n15012);
   U13221 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_5_port, B1 => 
                           n15145, B2 => REGISTERS_8_5_port, ZN => n15011);
   U13222 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_5_port, B1 => 
                           n15154, B2 => REGISTERS_21_5_port, ZN => n15010);
   U13223 : NAND4_X1 port map( A1 => n15013, A2 => n15012, A3 => n15011, A4 => 
                           n15010, ZN => n15014);
   U13224 : NOR3_X1 port map( A1 => n15016, A2 => n15015, A3 => n15014, ZN => 
                           n15017);
   U13225 : OAI222_X1 port map( A1 => n16026, A2 => n8447, B1 => n15115, B2 => 
                           n15018, C1 => n14354, C2 => n15017, ZN => n8564);
   U13226 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_4_port, B1 => 
                           n15088, B2 => REGISTERS_5_4_port, ZN => n15023);
   U13227 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_4_port, B1 => 
                           n15116, B2 => REGISTERS_0_4_port, ZN => n15022);
   U13228 : AOI22_X1 port map( A1 => n15121, A2 => REGISTERS_3_4_port, B1 => 
                           n15091, B2 => REGISTERS_7_4_port, ZN => n15021);
   U13229 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_4_port, B1 => 
                           n14483, B2 => REGISTERS_4_4_port, ZN => n15020);
   U13230 : AND4_X1 port map( A1 => n15023, A2 => n15022, A3 => n15021, A4 => 
                           n15020, ZN => n15042);
   U13231 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_4_port, B1 => 
                           n15096, B2 => REGISTERS_28_4_port, ZN => n15027);
   U13232 : AOI22_X1 port map( A1 => n15144, A2 => REGISTERS_9_4_port, B1 => 
                           n15126, B2 => REGISTERS_29_4_port, ZN => n15026);
   U13233 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_4_port, B1 => 
                           n15142, B2 => REGISTERS_14_4_port, ZN => n15025);
   U13234 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_4_port, B1 => 
                           n15127, B2 => REGISTERS_24_4_port, ZN => n15024);
   U13235 : NAND4_X1 port map( A1 => n15027, A2 => n15026, A3 => n15025, A4 => 
                           n15024, ZN => n15040);
   U13236 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_4_port, B1 => 
                           n15154, B2 => REGISTERS_21_4_port, ZN => n15031);
   U13237 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_4_port, B1 => 
                           n15128, B2 => REGISTERS_22_4_port, ZN => n15030);
   U13238 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_4_port, B1 => 
                           n15140, B2 => REGISTERS_12_4_port, ZN => n15029);
   U13239 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_4_port, B1 => 
                           n15150, B2 => REGISTERS_10_4_port, ZN => n15028);
   U13240 : NAND4_X1 port map( A1 => n15031, A2 => n15030, A3 => n15029, A4 => 
                           n15028, ZN => n15039);
   U13241 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_4_port, B1 => 
                           n15032, B2 => REGISTERS_30_4_port, ZN => n15037);
   U13242 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_4_port, B1 => 
                           n15130, B2 => REGISTERS_16_4_port, ZN => n15036);
   U13243 : AOI22_X1 port map( A1 => n15033, A2 => REGISTERS_26_4_port, B1 => 
                           n15153, B2 => REGISTERS_20_4_port, ZN => n15035);
   U13244 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_4_port, B1 => 
                           n15145, B2 => REGISTERS_8_4_port, ZN => n15034);
   U13245 : NAND4_X1 port map( A1 => n15037, A2 => n15036, A3 => n15035, A4 => 
                           n15034, ZN => n15038);
   U13246 : NOR3_X1 port map( A1 => n15040, A2 => n15039, A3 => n15038, ZN => 
                           n15041);
   U13247 : OAI222_X1 port map( A1 => n16071, A2 => n8446, B1 => n14505, B2 => 
                           n15042, C1 => n15166, C2 => n15041, ZN => n8565);
   U13248 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_3_port, B1 => 
                           n15090, B2 => REGISTERS_3_3_port, ZN => n15047);
   U13249 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_3_port, B1 => 
                           n15043, B2 => REGISTERS_6_3_port, ZN => n15046);
   U13250 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_3_port, B1 => 
                           n15089, B2 => REGISTERS_0_3_port, ZN => n15045);
   U13251 : AOI22_X1 port map( A1 => n14483, A2 => REGISTERS_4_3_port, B1 => 
                           n15091, B2 => REGISTERS_7_3_port, ZN => n15044);
   U13252 : AND4_X1 port map( A1 => n15047, A2 => n15046, A3 => n15045, A4 => 
                           n15044, ZN => n15064);
   U13253 : AOI22_X1 port map( A1 => n15152, A2 => REGISTERS_31_3_port, B1 => 
                           n15126, B2 => REGISTERS_29_3_port, ZN => n15051);
   U13254 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_3_port, B1 => 
                           n15156, B2 => REGISTERS_23_3_port, ZN => n15050);
   U13255 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_3_port, B1 => 
                           n15144, B2 => REGISTERS_9_3_port, ZN => n15049);
   U13256 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_3_port, B1 => 
                           n15128, B2 => REGISTERS_22_3_port, ZN => n15048);
   U13257 : NAND4_X1 port map( A1 => n15051, A2 => n15050, A3 => n15049, A4 => 
                           n15048, ZN => n15062);
   U13258 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_3_port, B1 => 
                           n15074, B2 => REGISTERS_30_3_port, ZN => n15055);
   U13259 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_3_port, B1 => 
                           n15150, B2 => REGISTERS_10_3_port, ZN => n15054);
   U13260 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_3_port, B1 => 
                           n15140, B2 => REGISTERS_12_3_port, ZN => n15053);
   U13261 : AOI22_X1 port map( A1 => n15151, A2 => REGISTERS_28_3_port, B1 => 
                           n15154, B2 => REGISTERS_21_3_port, ZN => n15052);
   U13262 : NAND4_X1 port map( A1 => n15055, A2 => n15054, A3 => n15053, A4 => 
                           n15052, ZN => n15061);
   U13263 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_3_port, B1 => 
                           n15143, B2 => REGISTERS_27_3_port, ZN => n15059);
   U13264 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_3_port, B1 => 
                           n15127, B2 => REGISTERS_24_3_port, ZN => n15058);
   U13265 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_3_port, B1 => 
                           n15145, B2 => REGISTERS_8_3_port, ZN => n15057);
   U13266 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_3_port, B1 => 
                           n15142, B2 => REGISTERS_14_3_port, ZN => n15056);
   U13267 : NAND4_X1 port map( A1 => n15059, A2 => n15058, A3 => n15057, A4 => 
                           n15056, ZN => n15060);
   U13268 : NOR3_X1 port map( A1 => n15062, A2 => n15061, A3 => n15060, ZN => 
                           n15063);
   U13269 : OAI222_X1 port map( A1 => n16026, A2 => n8445, B1 => n15115, B2 => 
                           n15064, C1 => n14354, C2 => n15063, ZN => n8566);
   U13270 : AOI22_X1 port map( A1 => n15088, A2 => REGISTERS_5_2_port, B1 => 
                           n15116, B2 => REGISTERS_0_2_port, ZN => n15069);
   U13271 : AOI22_X1 port map( A1 => n15090, A2 => REGISTERS_3_2_port, B1 => 
                           n15043, B2 => REGISTERS_6_2_port, ZN => n15068);
   U13272 : AOI22_X1 port map( A1 => n15065, A2 => REGISTERS_1_2_port, B1 => 
                           n14483, B2 => REGISTERS_4_2_port, ZN => n15067);
   U13273 : AOI22_X1 port map( A1 => n14506, A2 => REGISTERS_2_2_port, B1 => 
                           n15119, B2 => REGISTERS_7_2_port, ZN => n15066);
   U13274 : AND4_X1 port map( A1 => n15069, A2 => n15068, A3 => n15067, A4 => 
                           n15066, ZN => n15087);
   U13275 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_2_port, B1 => 
                           n15128, B2 => REGISTERS_22_2_port, ZN => n15073);
   U13276 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_2_port, B1 => 
                           n15096, B2 => REGISTERS_28_2_port, ZN => n15072);
   U13277 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_2_port, B1 => 
                           n15143, B2 => REGISTERS_27_2_port, ZN => n15071);
   U13278 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_2_port, B1 => 
                           n15142, B2 => REGISTERS_14_2_port, ZN => n15070);
   U13279 : NAND4_X1 port map( A1 => n15073, A2 => n15072, A3 => n15071, A4 => 
                           n15070, ZN => n15085);
   U13280 : AOI22_X1 port map( A1 => n15150, A2 => REGISTERS_10_2_port, B1 => 
                           n15144, B2 => REGISTERS_9_2_port, ZN => n15078);
   U13281 : AOI22_X1 port map( A1 => n15130, A2 => REGISTERS_16_2_port, B1 => 
                           n15145, B2 => REGISTERS_8_2_port, ZN => n15077);
   U13282 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_2_port, B1 => 
                           n15156, B2 => REGISTERS_23_2_port, ZN => n15076);
   U13283 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_2_port, B1 => 
                           n15074, B2 => REGISTERS_30_2_port, ZN => n15075);
   U13284 : NAND4_X1 port map( A1 => n15078, A2 => n15077, A3 => n15076, A4 => 
                           n15075, ZN => n15084);
   U13285 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_2_port, B1 => 
                           n15140, B2 => REGISTERS_12_2_port, ZN => n15082);
   U13286 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_2_port, B1 => 
                           n15152, B2 => REGISTERS_31_2_port, ZN => n15081);
   U13287 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_2_port, B1 => 
                           n15126, B2 => REGISTERS_29_2_port, ZN => n15080);
   U13288 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_2_port, B1 => 
                           n15154, B2 => REGISTERS_21_2_port, ZN => n15079);
   U13289 : NAND4_X1 port map( A1 => n15082, A2 => n15081, A3 => n15080, A4 => 
                           n15079, ZN => n15083);
   U13290 : NOR3_X1 port map( A1 => n15085, A2 => n15084, A3 => n15083, ZN => 
                           n15086);
   U13291 : OAI222_X1 port map( A1 => n16071, A2 => n8444, B1 => n15115, B2 => 
                           n15087, C1 => n15166, C2 => n15086, ZN => n8567);
   U13292 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_1_port, B1 => 
                           n15088, B2 => REGISTERS_5_1_port, ZN => n15095);
   U13293 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_1_port, B1 => 
                           n15089, B2 => REGISTERS_0_1_port, ZN => n15094);
   U13294 : AOI22_X1 port map( A1 => n15019, A2 => REGISTERS_2_1_port, B1 => 
                           n15090, B2 => REGISTERS_3_1_port, ZN => n15093);
   U13295 : AOI22_X1 port map( A1 => n14483, A2 => REGISTERS_4_1_port, B1 => 
                           n15091, B2 => REGISTERS_7_1_port, ZN => n15092);
   U13296 : AND4_X1 port map( A1 => n15095, A2 => n15094, A3 => n15093, A4 => 
                           n15092, ZN => n15114);
   U13297 : AOI22_X1 port map( A1 => n15156, A2 => REGISTERS_23_1_port, B1 => 
                           n15154, B2 => REGISTERS_21_1_port, ZN => n15100);
   U13298 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_1_port, B1 => 
                           n15096, B2 => REGISTERS_28_1_port, ZN => n15099);
   U13299 : AOI22_X1 port map( A1 => n15132, A2 => REGISTERS_15_1_port, B1 => 
                           n15130, B2 => REGISTERS_16_1_port, ZN => n15098);
   U13300 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_1_port, B1 => 
                           n15140, B2 => REGISTERS_12_1_port, ZN => n15097);
   U13301 : NAND4_X1 port map( A1 => n15100, A2 => n15099, A3 => n15098, A4 => 
                           n15097, ZN => n15112);
   U13302 : AOI22_X1 port map( A1 => n15138, A2 => REGISTERS_11_1_port, B1 => 
                           n15127, B2 => REGISTERS_24_1_port, ZN => n15105);
   U13303 : AOI22_X1 port map( A1 => n15101, A2 => REGISTERS_18_1_port, B1 => 
                           n15150, B2 => REGISTERS_10_1_port, ZN => n15104);
   U13304 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_1_port, B1 => 
                           n15128, B2 => REGISTERS_22_1_port, ZN => n15103);
   U13305 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_1_port, B1 => 
                           n15144, B2 => REGISTERS_9_1_port, ZN => n15102);
   U13306 : NAND4_X1 port map( A1 => n15105, A2 => n15104, A3 => n15103, A4 => 
                           n15102, ZN => n15111);
   U13307 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_1_port, B1 => 
                           n15145, B2 => REGISTERS_8_1_port, ZN => n15109);
   U13308 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_1_port, B1 => 
                           n15152, B2 => REGISTERS_31_1_port, ZN => n15108);
   U13309 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_1_port, B1 => 
                           n15142, B2 => REGISTERS_14_1_port, ZN => n15107);
   U13310 : AOI22_X1 port map( A1 => n14832, A2 => REGISTERS_19_1_port, B1 => 
                           n15126, B2 => REGISTERS_29_1_port, ZN => n15106);
   U13311 : NAND4_X1 port map( A1 => n15109, A2 => n15108, A3 => n15107, A4 => 
                           n15106, ZN => n15110);
   U13312 : NOR3_X1 port map( A1 => n15112, A2 => n15111, A3 => n15110, ZN => 
                           n15113);
   U13313 : OAI222_X1 port map( A1 => n16026, A2 => n8443, B1 => n15115, B2 => 
                           n15114, C1 => n14354, C2 => n15113, ZN => n8568);
   U13314 : AOI22_X1 port map( A1 => n15043, A2 => REGISTERS_6_0_port, B1 => 
                           n15116, B2 => REGISTERS_0_0_port, ZN => n15125);
   U13315 : AOI22_X1 port map( A1 => n15118, A2 => REGISTERS_5_0_port, B1 => 
                           n15117, B2 => REGISTERS_4_0_port, ZN => n15124);
   U13316 : AOI22_X1 port map( A1 => n15120, A2 => REGISTERS_1_0_port, B1 => 
                           n15119, B2 => REGISTERS_7_0_port, ZN => n15123);
   U13317 : AOI22_X1 port map( A1 => n14759, A2 => REGISTERS_2_0_port, B1 => 
                           n15121, B2 => REGISTERS_3_0_port, ZN => n15122);
   U13318 : AND4_X1 port map( A1 => n15125, A2 => n15124, A3 => n15123, A4 => 
                           n15122, ZN => n15167);
   U13319 : AOI22_X1 port map( A1 => n15127, A2 => REGISTERS_24_0_port, B1 => 
                           n15126, B2 => REGISTERS_29_0_port, ZN => n15137);
   U13320 : AOI22_X1 port map( A1 => n15129, A2 => REGISTERS_17_0_port, B1 => 
                           n15128, B2 => REGISTERS_22_0_port, ZN => n15136);
   U13321 : AOI22_X1 port map( A1 => n15131, A2 => REGISTERS_26_0_port, B1 => 
                           n15130, B2 => REGISTERS_16_0_port, ZN => n15135);
   U13322 : AOI22_X1 port map( A1 => n15133, A2 => REGISTERS_30_0_port, B1 => 
                           n15132, B2 => REGISTERS_15_0_port, ZN => n15134);
   U13323 : NAND4_X1 port map( A1 => n15137, A2 => n15136, A3 => n15135, A4 => 
                           n15134, ZN => n15164);
   U13324 : AOI22_X1 port map( A1 => n15139, A2 => REGISTERS_19_0_port, B1 => 
                           n15138, B2 => REGISTERS_11_0_port, ZN => n15149);
   U13325 : AOI22_X1 port map( A1 => n15141, A2 => REGISTERS_25_0_port, B1 => 
                           n15140, B2 => REGISTERS_12_0_port, ZN => n15148);
   U13326 : AOI22_X1 port map( A1 => n15143, A2 => REGISTERS_27_0_port, B1 => 
                           n15142, B2 => REGISTERS_14_0_port, ZN => n15147);
   U13327 : AOI22_X1 port map( A1 => n15145, A2 => REGISTERS_8_0_port, B1 => 
                           n15144, B2 => REGISTERS_9_0_port, ZN => n15146);
   U13328 : NAND4_X1 port map( A1 => n15149, A2 => n15148, A3 => n15147, A4 => 
                           n15146, ZN => n15163);
   U13329 : AOI22_X1 port map( A1 => n15151, A2 => REGISTERS_28_0_port, B1 => 
                           n15150, B2 => REGISTERS_10_0_port, ZN => n15161);
   U13330 : AOI22_X1 port map( A1 => n15153, A2 => REGISTERS_20_0_port, B1 => 
                           n15152, B2 => REGISTERS_31_0_port, ZN => n15160);
   U13331 : AOI22_X1 port map( A1 => n15155, A2 => REGISTERS_18_0_port, B1 => 
                           n15154, B2 => REGISTERS_21_0_port, ZN => n15159);
   U13332 : AOI22_X1 port map( A1 => n15157, A2 => REGISTERS_13_0_port, B1 => 
                           n15156, B2 => REGISTERS_23_0_port, ZN => n15158);
   U13333 : NAND4_X1 port map( A1 => n15161, A2 => n15160, A3 => n15159, A4 => 
                           n15158, ZN => n15162);
   U13334 : NOR3_X1 port map( A1 => n15164, A2 => n15163, A3 => n15162, ZN => 
                           n15165);
   U13335 : OAI222_X1 port map( A1 => n16071, A2 => n8442, B1 => n14505, B2 => 
                           n15167, C1 => n15166, C2 => n15165, ZN => n8569);
   U13336 : NAND3_X1 port map( A1 => ENABLE, A2 => RD2, A3 => n13731, ZN => 
                           n16605);
   U13337 : CLKBUF_X2 port map( A => n16605, Z => n15796);
   U13338 : INV_X1 port map( A => ADD_RD2(0), ZN => n15185);
   U13339 : INV_X1 port map( A => ADD_RD2(1), ZN => n15188);
   U13340 : NOR3_X1 port map( A1 => n15185, A2 => n15188, A3 => ADD_RD2(2), ZN 
                           => n15746);
   U13341 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => n15168, ZN => n15204);
   U13342 : NOR2_X1 port map( A1 => n15301, A2 => n15204, ZN => n16530);
   U13343 : CLKBUF_X2 port map( A => n16530, Z => n16414);
   U13344 : OR2_X1 port map( A1 => n15168, A2 => ADD_RD2(3), ZN => n15202);
   U13345 : NOR2_X1 port map( A1 => n15202, A2 => n15236, ZN => n15169);
   U13346 : AOI22_X1 port map( A1 => REGISTERS_11_63_port, A2 => n16414, B1 => 
                           REGISTERS_20_63_port, B2 => n16581, ZN => n15179);
   U13347 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n15199
                           );
   U13348 : NOR3_X1 port map( A1 => n15185, A2 => ADD_RD2(1), A3 => ADD_RD2(2),
                           ZN => n16322);
   U13349 : NOR2_X1 port map( A1 => n15199, A2 => n15556, ZN => n15170);
   U13350 : NOR3_X1 port map( A1 => n15188, A2 => n15184, A3 => ADD_RD2(0), ZN 
                           => n16344);
   U13351 : NOR2_X1 port map( A1 => n15199, A2 => n15258, ZN => n15171);
   U13352 : AOI22_X1 port map( A1 => REGISTERS_25_63_port, A2 => n16557, B1 => 
                           REGISTERS_30_63_port, B2 => n16555, ZN => n15178);
   U13353 : NOR2_X1 port map( A1 => n15202, A2 => n15556, ZN => n15172);
   U13354 : NOR2_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), ZN => n15189)
                           ;
   U13355 : NAND2_X1 port map( A1 => ADD_RD2(1), A2 => n15189, ZN => n15214);
   U13356 : NOR2_X1 port map( A1 => n15214, A2 => n15204, ZN => n15173);
   U13357 : AOI22_X1 port map( A1 => REGISTERS_17_63_port, A2 => n16579, B1 => 
                           REGISTERS_10_63_port, B2 => n16560, ZN => n15177);
   U13358 : NOR2_X1 port map( A1 => n15204, A2 => n15236, ZN => n15174);
   U13359 : NOR3_X1 port map( A1 => n15185, A2 => n15184, A3 => ADD_RD2(1), ZN 
                           => n16215);
   U13360 : NOR2_X1 port map( A1 => n15202, A2 => n15344, ZN => n15175);
   U13361 : AOI22_X1 port map( A1 => REGISTERS_12_63_port, A2 => n16580, B1 => 
                           REGISTERS_21_63_port, B2 => n16568, ZN => n15176);
   U13362 : NAND4_X1 port map( A1 => n15179, A2 => n15178, A3 => n15177, A4 => 
                           n15176, ZN => n15212);
   U13363 : NOR2_X1 port map( A1 => n15199, A2 => n15214, ZN => n15180);
   U13364 : NOR2_X1 port map( A1 => n15204, A2 => n15344, ZN => n15181);
   U13365 : AOI22_X1 port map( A1 => REGISTERS_26_63_port, A2 => n16582, B1 => 
                           REGISTERS_13_63_port, B2 => n16562, ZN => n15194);
   U13366 : NOR2_X1 port map( A1 => n15199, A2 => n15236, ZN => n15182);
   U13367 : NOR2_X1 port map( A1 => n15199, A2 => n15344, ZN => n15183);
   U13368 : AOI22_X1 port map( A1 => REGISTERS_28_63_port, A2 => n16570, B1 => 
                           REGISTERS_29_63_port, B2 => n16574, ZN => n15193);
   U13369 : NOR3_X1 port map( A1 => n15188, A2 => n15185, A3 => n15184, ZN => 
                           n16216);
   U13370 : NOR2_X1 port map( A1 => n15202, A2 => n15366, ZN => n15186);
   U13371 : NOR2_X1 port map( A1 => n15204, A2 => n15556, ZN => n16437);
   U13372 : CLKBUF_X2 port map( A => n16437, Z => n16029);
   U13373 : CLKBUF_X2 port map( A => n16029, Z => n16525);
   U13374 : AOI22_X1 port map( A1 => REGISTERS_23_63_port, A2 => n16572, B1 => 
                           REGISTERS_9_63_port, B2 => n16525, ZN => n15192);
   U13375 : NOR2_X1 port map( A1 => n15204, A2 => n15366, ZN => n15187);
   U13376 : NAND2_X1 port map( A1 => n15189, A2 => n15188, ZN => n15213);
   U13377 : NOR2_X1 port map( A1 => n15199, A2 => n15213, ZN => n15190);
   U13378 : AOI22_X1 port map( A1 => REGISTERS_15_63_port, A2 => n16558, B1 => 
                           REGISTERS_24_63_port, B2 => n16559, ZN => n15191);
   U13379 : NAND4_X1 port map( A1 => n15194, A2 => n15193, A3 => n15192, A4 => 
                           n15191, ZN => n15211);
   U13380 : NOR2_X1 port map( A1 => n15202, A2 => n15214, ZN => n15195);
   U13381 : NOR2_X1 port map( A1 => n15202, A2 => n15258, ZN => n15196);
   U13382 : AOI22_X1 port map( A1 => REGISTERS_18_63_port, A2 => n16584, B1 => 
                           REGISTERS_22_63_port, B2 => n16556, ZN => n15209);
   U13383 : NOR2_X1 port map( A1 => n15202, A2 => n15301, ZN => n15197);
   U13384 : NOR2_X1 port map( A1 => n15301, A2 => n15199, ZN => n15198);
   U13385 : AOI22_X1 port map( A1 => REGISTERS_19_63_port, A2 => n16569, B1 => 
                           REGISTERS_27_63_port, B2 => n16573, ZN => n15208);
   U13386 : NOR2_X1 port map( A1 => n15199, A2 => n15366, ZN => n15200);
   U13387 : NOR2_X1 port map( A1 => n15213, A2 => n15204, ZN => n15201);
   U13388 : AOI22_X1 port map( A1 => REGISTERS_31_63_port, A2 => n16583, B1 => 
                           REGISTERS_8_63_port, B2 => n16567, ZN => n15207);
   U13389 : NOR2_X1 port map( A1 => n15202, A2 => n15213, ZN => n15203);
   U13390 : NOR2_X1 port map( A1 => n15258, A2 => n15204, ZN => n15205);
   U13391 : AOI22_X1 port map( A1 => REGISTERS_16_63_port, A2 => n16561, B1 => 
                           REGISTERS_14_63_port, B2 => n16571, ZN => n15206);
   U13392 : NAND4_X1 port map( A1 => n15209, A2 => n15208, A3 => n15207, A4 => 
                           n15206, ZN => n15210);
   U13393 : NOR3_X1 port map( A1 => n15212, A2 => n15211, A3 => n15210, ZN => 
                           n15220);
   U13394 : OR3_X2 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n16605, 
                           ZN => n16553);
   U13395 : INV_X2 port map( A => n15556, ZN => n16544);
   U13396 : INV_X2 port map( A => n15213, ZN => n16547);
   U13397 : AOI22_X1 port map( A1 => REGISTERS_1_63_port, A2 => n16544, B1 => 
                           REGISTERS_0_63_port, B2 => n16597, ZN => n15218);
   U13398 : INV_X2 port map( A => n15344, ZN => n16518);
   U13399 : AOI22_X1 port map( A1 => REGISTERS_3_63_port, A2 => n15746, B1 => 
                           REGISTERS_5_63_port, B2 => n16518, ZN => n15217);
   U13400 : INV_X2 port map( A => n15366, ZN => n16454);
   U13401 : AOI22_X1 port map( A1 => REGISTERS_7_63_port, A2 => n16454, B1 => 
                           REGISTERS_6_63_port, B2 => n16592, ZN => n15216);
   U13402 : INV_X2 port map( A => n15214, ZN => n16545);
   U13403 : INV_X2 port map( A => n15236, ZN => n16543);
   U13404 : AOI22_X1 port map( A1 => REGISTERS_2_63_port, A2 => n16545, B1 => 
                           REGISTERS_4_63_port, B2 => n16543, ZN => n15215);
   U13405 : OAI222_X1 port map( A1 => n15796, A2 => n15220, B1 => n16553, B2 =>
                           n15219, C1 => n14910, C2 => n8441, ZN => n8570);
   U13406 : AOI22_X1 port map( A1 => REGISTERS_8_62_port, A2 => n16567, B1 => 
                           REGISTERS_12_62_port, B2 => n16580, ZN => n15224);
   U13407 : AOI22_X1 port map( A1 => REGISTERS_24_62_port, A2 => n16559, B1 => 
                           REGISTERS_22_62_port, B2 => n16556, ZN => n15223);
   U13408 : AOI22_X1 port map( A1 => REGISTERS_17_62_port, A2 => n16579, B1 => 
                           REGISTERS_31_62_port, B2 => n16583, ZN => n15222);
   U13409 : AOI22_X1 port map( A1 => REGISTERS_27_62_port, A2 => n16573, B1 => 
                           REGISTERS_23_62_port, B2 => n16572, ZN => n15221);
   U13410 : NAND4_X1 port map( A1 => n15224, A2 => n15223, A3 => n15222, A4 => 
                           n15221, ZN => n15235);
   U13411 : AOI22_X1 port map( A1 => REGISTERS_13_62_port, A2 => n16562, B1 => 
                           REGISTERS_20_62_port, B2 => n16581, ZN => n15228);
   U13412 : AOI22_X1 port map( A1 => REGISTERS_11_62_port, A2 => n16530, B1 => 
                           REGISTERS_9_62_port, B2 => n16525, ZN => n15227);
   U13413 : AOI22_X1 port map( A1 => REGISTERS_16_62_port, A2 => n16561, B1 => 
                           REGISTERS_21_62_port, B2 => n16568, ZN => n15226);
   U13414 : AOI22_X1 port map( A1 => REGISTERS_26_62_port, A2 => n16582, B1 => 
                           REGISTERS_25_62_port, B2 => n16557, ZN => n15225);
   U13415 : NAND4_X1 port map( A1 => n15228, A2 => n15227, A3 => n15226, A4 => 
                           n15225, ZN => n15234);
   U13416 : AOI22_X1 port map( A1 => REGISTERS_29_62_port, A2 => n16574, B1 => 
                           REGISTERS_19_62_port, B2 => n16569, ZN => n15232);
   U13417 : AOI22_X1 port map( A1 => REGISTERS_18_62_port, A2 => n16584, B1 => 
                           REGISTERS_30_62_port, B2 => n16555, ZN => n15231);
   U13418 : AOI22_X1 port map( A1 => REGISTERS_10_62_port, A2 => n16560, B1 => 
                           REGISTERS_14_62_port, B2 => n16571, ZN => n15230);
   U13419 : AOI22_X1 port map( A1 => REGISTERS_15_62_port, A2 => n16558, B1 => 
                           REGISTERS_28_62_port, B2 => n16570, ZN => n15229);
   U13420 : NAND4_X1 port map( A1 => n15232, A2 => n15231, A3 => n15230, A4 => 
                           n15229, ZN => n15233);
   U13421 : NOR3_X1 port map( A1 => n15235, A2 => n15234, A3 => n15233, ZN => 
                           n15242);
   U13422 : INV_X2 port map( A => n15258, ZN => n16546);
   U13423 : AOI22_X1 port map( A1 => REGISTERS_2_62_port, A2 => n16596, B1 => 
                           REGISTERS_6_62_port, B2 => n16546, ZN => n15240);
   U13424 : AOI22_X1 port map( A1 => REGISTERS_4_62_port, A2 => n16543, B1 => 
                           REGISTERS_0_62_port, B2 => n16547, ZN => n15239);
   U13425 : INV_X2 port map( A => n15301, ZN => n16453);
   U13426 : AOI22_X1 port map( A1 => REGISTERS_3_62_port, A2 => n16453, B1 => 
                           REGISTERS_5_62_port, B2 => n16518, ZN => n15238);
   U13427 : AOI22_X1 port map( A1 => REGISTERS_7_62_port, A2 => n16454, B1 => 
                           REGISTERS_1_62_port, B2 => n16430, ZN => n15237);
   U13428 : AND4_X1 port map( A1 => n15240, A2 => n15239, A3 => n15238, A4 => 
                           n15237, ZN => n15241);
   U13429 : OAI222_X1 port map( A1 => n16605, A2 => n15242, B1 => n16603, B2 =>
                           n15241, C1 => n16071, C2 => n8440, ZN => n8571);
   U13430 : AOI22_X1 port map( A1 => REGISTERS_14_61_port, A2 => n16571, B1 => 
                           REGISTERS_26_61_port, B2 => n16582, ZN => n15246);
   U13431 : AOI22_X1 port map( A1 => REGISTERS_16_61_port, A2 => n16561, B1 => 
                           REGISTERS_28_61_port, B2 => n16570, ZN => n15245);
   U13432 : AOI22_X1 port map( A1 => REGISTERS_21_61_port, A2 => n16568, B1 => 
                           REGISTERS_22_61_port, B2 => n16556, ZN => n15244);
   U13433 : AOI22_X1 port map( A1 => REGISTERS_29_61_port, A2 => n16574, B1 => 
                           REGISTERS_25_61_port, B2 => n16557, ZN => n15243);
   U13434 : NAND4_X1 port map( A1 => n15246, A2 => n15245, A3 => n15244, A4 => 
                           n15243, ZN => n15257);
   U13435 : AOI22_X1 port map( A1 => REGISTERS_9_61_port, A2 => n16437, B1 => 
                           REGISTERS_20_61_port, B2 => n16581, ZN => n15250);
   U13436 : AOI22_X1 port map( A1 => REGISTERS_8_61_port, A2 => n16567, B1 => 
                           REGISTERS_10_61_port, B2 => n16560, ZN => n15249);
   U13437 : AOI22_X1 port map( A1 => REGISTERS_13_61_port, A2 => n16562, B1 => 
                           REGISTERS_18_61_port, B2 => n16584, ZN => n15248);
   U13438 : AOI22_X1 port map( A1 => REGISTERS_15_61_port, A2 => n16558, B1 => 
                           REGISTERS_30_61_port, B2 => n16555, ZN => n15247);
   U13439 : NAND4_X1 port map( A1 => n15250, A2 => n15249, A3 => n15248, A4 => 
                           n15247, ZN => n15256);
   U13440 : AOI22_X1 port map( A1 => REGISTERS_19_61_port, A2 => n16569, B1 => 
                           REGISTERS_27_61_port, B2 => n16573, ZN => n15254);
   U13441 : AOI22_X1 port map( A1 => REGISTERS_24_61_port, A2 => n16559, B1 => 
                           REGISTERS_12_61_port, B2 => n16580, ZN => n15253);
   U13442 : AOI22_X1 port map( A1 => REGISTERS_11_61_port, A2 => n16530, B1 => 
                           REGISTERS_17_61_port, B2 => n16579, ZN => n15252);
   U13443 : AOI22_X1 port map( A1 => REGISTERS_23_61_port, A2 => n16572, B1 => 
                           REGISTERS_31_61_port, B2 => n16583, ZN => n15251);
   U13444 : NAND4_X1 port map( A1 => n15254, A2 => n15253, A3 => n15252, A4 => 
                           n15251, ZN => n15255);
   U13445 : NOR3_X1 port map( A1 => n15257, A2 => n15256, A3 => n15255, ZN => 
                           n15264);
   U13446 : AOI22_X1 port map( A1 => REGISTERS_7_61_port, A2 => n16454, B1 => 
                           REGISTERS_5_61_port, B2 => n16518, ZN => n15262);
   U13447 : AOI22_X1 port map( A1 => REGISTERS_1_61_port, A2 => n16544, B1 => 
                           REGISTERS_4_61_port, B2 => n16543, ZN => n15261);
   U13448 : AOI22_X1 port map( A1 => REGISTERS_6_61_port, A2 => n16592, B1 => 
                           REGISTERS_3_61_port, B2 => n16593, ZN => n15260);
   U13449 : AOI22_X1 port map( A1 => REGISTERS_0_61_port, A2 => n16547, B1 => 
                           REGISTERS_2_61_port, B2 => n16596, ZN => n15259);
   U13450 : AND4_X1 port map( A1 => n15262, A2 => n15261, A3 => n15260, A4 => 
                           n15259, ZN => n15263);
   U13451 : OAI222_X1 port map( A1 => n15796, A2 => n15264, B1 => n16553, B2 =>
                           n15263, C1 => n16071, C2 => n8439, ZN => n8572);
   U13452 : AOI22_X1 port map( A1 => REGISTERS_12_60_port, A2 => n16580, B1 => 
                           REGISTERS_17_60_port, B2 => n16579, ZN => n15268);
   U13453 : AOI22_X1 port map( A1 => REGISTERS_19_60_port, A2 => n16569, B1 => 
                           REGISTERS_28_60_port, B2 => n16570, ZN => n15267);
   U13454 : AOI22_X1 port map( A1 => REGISTERS_13_60_port, A2 => n16562, B1 => 
                           REGISTERS_20_60_port, B2 => n16581, ZN => n15266);
   U13455 : AOI22_X1 port map( A1 => REGISTERS_24_60_port, A2 => n16559, B1 => 
                           REGISTERS_16_60_port, B2 => n16561, ZN => n15265);
   U13456 : NAND4_X1 port map( A1 => n15268, A2 => n15267, A3 => n15266, A4 => 
                           n15265, ZN => n15279);
   U13457 : AOI22_X1 port map( A1 => REGISTERS_30_60_port, A2 => n16555, B1 => 
                           REGISTERS_10_60_port, B2 => n16560, ZN => n15272);
   U13458 : AOI22_X1 port map( A1 => REGISTERS_14_60_port, A2 => n16571, B1 => 
                           REGISTERS_23_60_port, B2 => n16572, ZN => n15271);
   U13459 : AOI22_X1 port map( A1 => REGISTERS_29_60_port, A2 => n16574, B1 => 
                           REGISTERS_18_60_port, B2 => n16584, ZN => n15270);
   U13460 : AOI22_X1 port map( A1 => REGISTERS_22_60_port, A2 => n16556, B1 => 
                           REGISTERS_21_60_port, B2 => n16568, ZN => n15269);
   U13461 : NAND4_X1 port map( A1 => n15272, A2 => n15271, A3 => n15270, A4 => 
                           n15269, ZN => n15278);
   U13462 : AOI22_X1 port map( A1 => REGISTERS_9_60_port, A2 => n16437, B1 => 
                           REGISTERS_31_60_port, B2 => n16583, ZN => n15276);
   U13463 : CLKBUF_X2 port map( A => n16530, Z => n15782);
   U13464 : AOI22_X1 port map( A1 => REGISTERS_8_60_port, A2 => n16567, B1 => 
                           REGISTERS_11_60_port, B2 => n15782, ZN => n15275);
   U13465 : AOI22_X1 port map( A1 => REGISTERS_15_60_port, A2 => n16558, B1 => 
                           REGISTERS_26_60_port, B2 => n16582, ZN => n15274);
   U13466 : AOI22_X1 port map( A1 => REGISTERS_25_60_port, A2 => n16557, B1 => 
                           REGISTERS_27_60_port, B2 => n16573, ZN => n15273);
   U13467 : NAND4_X1 port map( A1 => n15276, A2 => n15275, A3 => n15274, A4 => 
                           n15273, ZN => n15277);
   U13468 : NOR3_X1 port map( A1 => n15279, A2 => n15278, A3 => n15277, ZN => 
                           n15285);
   U13469 : AOI22_X1 port map( A1 => REGISTERS_3_60_port, A2 => n16453, B1 => 
                           REGISTERS_6_60_port, B2 => n16546, ZN => n15283);
   U13470 : AOI22_X1 port map( A1 => REGISTERS_2_60_port, A2 => n16545, B1 => 
                           REGISTERS_5_60_port, B2 => n16518, ZN => n15282);
   U13471 : AOI22_X1 port map( A1 => REGISTERS_4_60_port, A2 => n16595, B1 => 
                           REGISTERS_0_60_port, B2 => n16547, ZN => n15281);
   U13472 : AOI22_X1 port map( A1 => REGISTERS_7_60_port, A2 => n16454, B1 => 
                           REGISTERS_1_60_port, B2 => n16544, ZN => n15280);
   U13473 : AND4_X1 port map( A1 => n15283, A2 => n15282, A3 => n15281, A4 => 
                           n15280, ZN => n15284);
   U13474 : OAI222_X1 port map( A1 => n16605, A2 => n15285, B1 => n16603, B2 =>
                           n15284, C1 => n16026, C2 => n8438, ZN => n8573);
   U13475 : AOI22_X1 port map( A1 => REGISTERS_25_59_port, A2 => n16557, B1 => 
                           REGISTERS_15_59_port, B2 => n16558, ZN => n15289);
   U13476 : AOI22_X1 port map( A1 => REGISTERS_11_59_port, A2 => n16414, B1 => 
                           REGISTERS_20_59_port, B2 => n16581, ZN => n15288);
   U13477 : AOI22_X1 port map( A1 => REGISTERS_24_59_port, A2 => n16559, B1 => 
                           REGISTERS_19_59_port, B2 => n16569, ZN => n15287);
   U13478 : AOI22_X1 port map( A1 => REGISTERS_13_59_port, A2 => n16562, B1 => 
                           REGISTERS_10_59_port, B2 => n16560, ZN => n15286);
   U13479 : NAND4_X1 port map( A1 => n15289, A2 => n15288, A3 => n15287, A4 => 
                           n15286, ZN => n15300);
   U13480 : AOI22_X1 port map( A1 => REGISTERS_27_59_port, A2 => n16573, B1 => 
                           REGISTERS_9_59_port, B2 => n16029, ZN => n15293);
   U13481 : AOI22_X1 port map( A1 => REGISTERS_26_59_port, A2 => n16582, B1 => 
                           REGISTERS_16_59_port, B2 => n16561, ZN => n15292);
   U13482 : AOI22_X1 port map( A1 => REGISTERS_14_59_port, A2 => n16571, B1 => 
                           REGISTERS_18_59_port, B2 => n16584, ZN => n15291);
   U13483 : AOI22_X1 port map( A1 => REGISTERS_22_59_port, A2 => n16556, B1 => 
                           REGISTERS_30_59_port, B2 => n16555, ZN => n15290);
   U13484 : NAND4_X1 port map( A1 => n15293, A2 => n15292, A3 => n15291, A4 => 
                           n15290, ZN => n15299);
   U13485 : AOI22_X1 port map( A1 => REGISTERS_31_59_port, A2 => n16583, B1 => 
                           REGISTERS_29_59_port, B2 => n16574, ZN => n15297);
   U13486 : AOI22_X1 port map( A1 => REGISTERS_28_59_port, A2 => n16570, B1 => 
                           REGISTERS_23_59_port, B2 => n16572, ZN => n15296);
   U13487 : AOI22_X1 port map( A1 => REGISTERS_21_59_port, A2 => n16568, B1 => 
                           REGISTERS_8_59_port, B2 => n16567, ZN => n15295);
   U13488 : AOI22_X1 port map( A1 => REGISTERS_12_59_port, A2 => n16580, B1 => 
                           REGISTERS_17_59_port, B2 => n16579, ZN => n15294);
   U13489 : NAND4_X1 port map( A1 => n15297, A2 => n15296, A3 => n15295, A4 => 
                           n15294, ZN => n15298);
   U13490 : NOR3_X1 port map( A1 => n15300, A2 => n15299, A3 => n15298, ZN => 
                           n15307);
   U13491 : AOI22_X1 port map( A1 => REGISTERS_1_59_port, A2 => n16544, B1 => 
                           REGISTERS_4_59_port, B2 => n16543, ZN => n15305);
   U13492 : AOI22_X1 port map( A1 => REGISTERS_0_59_port, A2 => n16597, B1 => 
                           REGISTERS_3_59_port, B2 => n16453, ZN => n15304);
   U13493 : AOI22_X1 port map( A1 => REGISTERS_2_59_port, A2 => n16596, B1 => 
                           REGISTERS_5_59_port, B2 => n16518, ZN => n15303);
   U13494 : AOI22_X1 port map( A1 => REGISTERS_6_59_port, A2 => n16546, B1 => 
                           REGISTERS_7_59_port, B2 => n16594, ZN => n15302);
   U13495 : AND4_X1 port map( A1 => n15305, A2 => n15304, A3 => n15303, A4 => 
                           n15302, ZN => n15306);
   U13496 : CLKBUF_X2 port map( A => n16049, Z => n16026);
   U13497 : OAI222_X1 port map( A1 => n15796, A2 => n15307, B1 => n16553, B2 =>
                           n15306, C1 => n16026, C2 => n8437, ZN => n8574);
   U13498 : AOI22_X1 port map( A1 => REGISTERS_14_58_port, A2 => n16571, B1 => 
                           REGISTERS_10_58_port, B2 => n16560, ZN => n15311);
   U13499 : AOI22_X1 port map( A1 => REGISTERS_21_58_port, A2 => n16568, B1 => 
                           REGISTERS_31_58_port, B2 => n16583, ZN => n15310);
   U13500 : AOI22_X1 port map( A1 => REGISTERS_25_58_port, A2 => n16557, B1 => 
                           REGISTERS_24_58_port, B2 => n16559, ZN => n15309);
   U13501 : AOI22_X1 port map( A1 => REGISTERS_15_58_port, A2 => n16558, B1 => 
                           REGISTERS_11_58_port, B2 => n16414, ZN => n15308);
   U13502 : NAND4_X1 port map( A1 => n15311, A2 => n15310, A3 => n15309, A4 => 
                           n15308, ZN => n15322);
   U13503 : AOI22_X1 port map( A1 => REGISTERS_20_58_port, A2 => n16581, B1 => 
                           REGISTERS_17_58_port, B2 => n16579, ZN => n15315);
   U13504 : AOI22_X1 port map( A1 => REGISTERS_13_58_port, A2 => n16562, B1 => 
                           REGISTERS_27_58_port, B2 => n16573, ZN => n15314);
   U13505 : AOI22_X1 port map( A1 => REGISTERS_8_58_port, A2 => n16567, B1 => 
                           REGISTERS_18_58_port, B2 => n16584, ZN => n15313);
   U13506 : AOI22_X1 port map( A1 => REGISTERS_19_58_port, A2 => n16569, B1 => 
                           REGISTERS_26_58_port, B2 => n16582, ZN => n15312);
   U13507 : NAND4_X1 port map( A1 => n15315, A2 => n15314, A3 => n15313, A4 => 
                           n15312, ZN => n15321);
   U13508 : AOI22_X1 port map( A1 => REGISTERS_28_58_port, A2 => n16570, B1 => 
                           REGISTERS_12_58_port, B2 => n16580, ZN => n15319);
   U13509 : AOI22_X1 port map( A1 => REGISTERS_23_58_port, A2 => n16572, B1 => 
                           REGISTERS_16_58_port, B2 => n16561, ZN => n15318);
   U13510 : AOI22_X1 port map( A1 => REGISTERS_22_58_port, A2 => n16556, B1 => 
                           REGISTERS_9_58_port, B2 => n16525, ZN => n15317);
   U13511 : AOI22_X1 port map( A1 => REGISTERS_30_58_port, A2 => n16555, B1 => 
                           REGISTERS_29_58_port, B2 => n16574, ZN => n15316);
   U13512 : NAND4_X1 port map( A1 => n15319, A2 => n15318, A3 => n15317, A4 => 
                           n15316, ZN => n15320);
   U13513 : NOR3_X1 port map( A1 => n15322, A2 => n15321, A3 => n15320, ZN => 
                           n15328);
   U13514 : AOI22_X1 port map( A1 => REGISTERS_2_58_port, A2 => n16596, B1 => 
                           REGISTERS_1_58_port, B2 => n16430, ZN => n15326);
   U13515 : AOI22_X1 port map( A1 => REGISTERS_5_58_port, A2 => n16542, B1 => 
                           REGISTERS_4_58_port, B2 => n16543, ZN => n15325);
   U13516 : AOI22_X1 port map( A1 => REGISTERS_6_58_port, A2 => n16546, B1 => 
                           REGISTERS_0_58_port, B2 => n16547, ZN => n15324);
   U13517 : AOI22_X1 port map( A1 => REGISTERS_3_58_port, A2 => n16453, B1 => 
                           REGISTERS_7_58_port, B2 => n16454, ZN => n15323);
   U13518 : AND4_X1 port map( A1 => n15326, A2 => n15325, A3 => n15324, A4 => 
                           n15323, ZN => n15327);
   U13519 : OAI222_X1 port map( A1 => n15796, A2 => n15328, B1 => n16603, B2 =>
                           n15327, C1 => n16026, C2 => n8436, ZN => n8575);
   U13520 : AOI22_X1 port map( A1 => REGISTERS_30_57_port, A2 => n16555, B1 => 
                           REGISTERS_15_57_port, B2 => n16558, ZN => n15332);
   U13521 : AOI22_X1 port map( A1 => REGISTERS_19_57_port, A2 => n16569, B1 => 
                           REGISTERS_29_57_port, B2 => n16574, ZN => n15331);
   U13522 : AOI22_X1 port map( A1 => REGISTERS_18_57_port, A2 => n16584, B1 => 
                           REGISTERS_25_57_port, B2 => n16557, ZN => n15330);
   U13523 : AOI22_X1 port map( A1 => REGISTERS_8_57_port, A2 => n16567, B1 => 
                           REGISTERS_27_57_port, B2 => n16573, ZN => n15329);
   U13524 : NAND4_X1 port map( A1 => n15332, A2 => n15331, A3 => n15330, A4 => 
                           n15329, ZN => n15343);
   U13525 : AOI22_X1 port map( A1 => REGISTERS_28_57_port, A2 => n16570, B1 => 
                           REGISTERS_14_57_port, B2 => n16571, ZN => n15336);
   U13526 : AOI22_X1 port map( A1 => REGISTERS_24_57_port, A2 => n16559, B1 => 
                           REGISTERS_26_57_port, B2 => n16582, ZN => n15335);
   U13527 : AOI22_X1 port map( A1 => REGISTERS_9_57_port, A2 => n16437, B1 => 
                           REGISTERS_10_57_port, B2 => n16560, ZN => n15334);
   U13528 : AOI22_X1 port map( A1 => REGISTERS_23_57_port, A2 => n16572, B1 => 
                           REGISTERS_11_57_port, B2 => n16414, ZN => n15333);
   U13529 : NAND4_X1 port map( A1 => n15336, A2 => n15335, A3 => n15334, A4 => 
                           n15333, ZN => n15342);
   U13530 : AOI22_X1 port map( A1 => REGISTERS_22_57_port, A2 => n16556, B1 => 
                           REGISTERS_13_57_port, B2 => n16562, ZN => n15340);
   U13531 : AOI22_X1 port map( A1 => REGISTERS_21_57_port, A2 => n16568, B1 => 
                           REGISTERS_12_57_port, B2 => n16580, ZN => n15339);
   U13532 : AOI22_X1 port map( A1 => REGISTERS_20_57_port, A2 => n16581, B1 => 
                           REGISTERS_16_57_port, B2 => n16561, ZN => n15338);
   U13533 : AOI22_X1 port map( A1 => REGISTERS_17_57_port, A2 => n16579, B1 => 
                           REGISTERS_31_57_port, B2 => n16583, ZN => n15337);
   U13534 : NAND4_X1 port map( A1 => n15340, A2 => n15339, A3 => n15338, A4 => 
                           n15337, ZN => n15341);
   U13535 : NOR3_X1 port map( A1 => n15343, A2 => n15342, A3 => n15341, ZN => 
                           n15350);
   U13536 : AOI22_X1 port map( A1 => REGISTERS_6_57_port, A2 => n16592, B1 => 
                           REGISTERS_0_57_port, B2 => n16547, ZN => n15348);
   U13537 : AOI22_X1 port map( A1 => REGISTERS_7_57_port, A2 => n16454, B1 => 
                           REGISTERS_5_57_port, B2 => n16518, ZN => n15347);
   U13538 : INV_X2 port map( A => n15236, ZN => n16595);
   U13539 : AOI22_X1 port map( A1 => REGISTERS_4_57_port, A2 => n16595, B1 => 
                           REGISTERS_2_57_port, B2 => n16596, ZN => n15346);
   U13540 : AOI22_X1 port map( A1 => REGISTERS_1_57_port, A2 => n16544, B1 => 
                           REGISTERS_3_57_port, B2 => n16593, ZN => n15345);
   U13541 : OAI222_X1 port map( A1 => n16605, A2 => n15350, B1 => n16553, B2 =>
                           n15349, C1 => n16049, C2 => n8435, ZN => n8576);
   U13542 : AOI22_X1 port map( A1 => REGISTERS_8_56_port, A2 => n16567, B1 => 
                           REGISTERS_23_56_port, B2 => n16572, ZN => n15354);
   U13543 : AOI22_X1 port map( A1 => REGISTERS_13_56_port, A2 => n16562, B1 => 
                           REGISTERS_10_56_port, B2 => n16560, ZN => n15353);
   U13544 : AOI22_X1 port map( A1 => REGISTERS_27_56_port, A2 => n16573, B1 => 
                           REGISTERS_30_56_port, B2 => n16555, ZN => n15352);
   U13545 : AOI22_X1 port map( A1 => REGISTERS_19_56_port, A2 => n16569, B1 => 
                           REGISTERS_15_56_port, B2 => n16558, ZN => n15351);
   U13546 : NAND4_X1 port map( A1 => n15354, A2 => n15353, A3 => n15352, A4 => 
                           n15351, ZN => n15365);
   U13547 : AOI22_X1 port map( A1 => REGISTERS_11_56_port, A2 => n16414, B1 => 
                           REGISTERS_25_56_port, B2 => n16557, ZN => n15358);
   U13548 : AOI22_X1 port map( A1 => REGISTERS_22_56_port, A2 => n16556, B1 => 
                           REGISTERS_12_56_port, B2 => n16580, ZN => n15357);
   U13549 : AOI22_X1 port map( A1 => REGISTERS_28_56_port, A2 => n16570, B1 => 
                           REGISTERS_29_56_port, B2 => n16574, ZN => n15356);
   U13550 : AOI22_X1 port map( A1 => REGISTERS_17_56_port, A2 => n16579, B1 => 
                           REGISTERS_20_56_port, B2 => n16581, ZN => n15355);
   U13551 : NAND4_X1 port map( A1 => n15358, A2 => n15357, A3 => n15356, A4 => 
                           n15355, ZN => n15364);
   U13552 : AOI22_X1 port map( A1 => REGISTERS_21_56_port, A2 => n16568, B1 => 
                           REGISTERS_24_56_port, B2 => n16559, ZN => n15362);
   U13553 : AOI22_X1 port map( A1 => REGISTERS_26_56_port, A2 => n16582, B1 => 
                           REGISTERS_9_56_port, B2 => n16029, ZN => n15361);
   U13554 : AOI22_X1 port map( A1 => REGISTERS_16_56_port, A2 => n16561, B1 => 
                           REGISTERS_18_56_port, B2 => n16584, ZN => n15360);
   U13555 : AOI22_X1 port map( A1 => REGISTERS_31_56_port, A2 => n16583, B1 => 
                           REGISTERS_14_56_port, B2 => n16571, ZN => n15359);
   U13556 : NAND4_X1 port map( A1 => n15362, A2 => n15361, A3 => n15360, A4 => 
                           n15359, ZN => n15363);
   U13557 : NOR3_X1 port map( A1 => n15365, A2 => n15364, A3 => n15363, ZN => 
                           n15372);
   U13558 : AOI22_X1 port map( A1 => REGISTERS_0_56_port, A2 => n16547, B1 => 
                           REGISTERS_4_56_port, B2 => n16543, ZN => n15370);
   U13559 : AOI22_X1 port map( A1 => REGISTERS_5_56_port, A2 => n16542, B1 => 
                           REGISTERS_2_56_port, B2 => n16545, ZN => n15369);
   U13560 : AOI22_X1 port map( A1 => REGISTERS_7_56_port, A2 => n16594, B1 => 
                           REGISTERS_3_56_port, B2 => n16593, ZN => n15368);
   U13561 : AOI22_X1 port map( A1 => REGISTERS_6_56_port, A2 => n16546, B1 => 
                           REGISTERS_1_56_port, B2 => n16544, ZN => n15367);
   U13562 : AND4_X1 port map( A1 => n15370, A2 => n15369, A3 => n15368, A4 => 
                           n15367, ZN => n15371);
   U13563 : OAI222_X1 port map( A1 => n15796, A2 => n15372, B1 => n16603, B2 =>
                           n15371, C1 => n16026, C2 => n8434, ZN => n8577);
   U13564 : AOI22_X1 port map( A1 => REGISTERS_10_55_port, A2 => n16560, B1 => 
                           REGISTERS_12_55_port, B2 => n16580, ZN => n15376);
   U13565 : AOI22_X1 port map( A1 => REGISTERS_26_55_port, A2 => n16582, B1 => 
                           REGISTERS_14_55_port, B2 => n16571, ZN => n15375);
   U13566 : AOI22_X1 port map( A1 => REGISTERS_9_55_port, A2 => n16029, B1 => 
                           REGISTERS_13_55_port, B2 => n16562, ZN => n15374);
   U13567 : AOI22_X1 port map( A1 => REGISTERS_11_55_port, A2 => n16530, B1 => 
                           REGISTERS_27_55_port, B2 => n16573, ZN => n15373);
   U13568 : NAND4_X1 port map( A1 => n15376, A2 => n15375, A3 => n15374, A4 => 
                           n15373, ZN => n15387);
   U13569 : AOI22_X1 port map( A1 => REGISTERS_25_55_port, A2 => n16557, B1 => 
                           REGISTERS_30_55_port, B2 => n16555, ZN => n15380);
   U13570 : AOI22_X1 port map( A1 => REGISTERS_31_55_port, A2 => n16583, B1 => 
                           REGISTERS_29_55_port, B2 => n16574, ZN => n15379);
   U13571 : AOI22_X1 port map( A1 => REGISTERS_21_55_port, A2 => n16568, B1 => 
                           REGISTERS_20_55_port, B2 => n16581, ZN => n15378);
   U13572 : AOI22_X1 port map( A1 => REGISTERS_24_55_port, A2 => n16559, B1 => 
                           REGISTERS_17_55_port, B2 => n16579, ZN => n15377);
   U13573 : NAND4_X1 port map( A1 => n15380, A2 => n15379, A3 => n15378, A4 => 
                           n15377, ZN => n15386);
   U13574 : AOI22_X1 port map( A1 => REGISTERS_18_55_port, A2 => n16584, B1 => 
                           REGISTERS_28_55_port, B2 => n16570, ZN => n15384);
   U13575 : AOI22_X1 port map( A1 => REGISTERS_16_55_port, A2 => n16561, B1 => 
                           REGISTERS_8_55_port, B2 => n16567, ZN => n15383);
   U13576 : AOI22_X1 port map( A1 => REGISTERS_22_55_port, A2 => n16556, B1 => 
                           REGISTERS_19_55_port, B2 => n16569, ZN => n15382);
   U13577 : AOI22_X1 port map( A1 => REGISTERS_15_55_port, A2 => n16558, B1 => 
                           REGISTERS_23_55_port, B2 => n16572, ZN => n15381);
   U13578 : NAND4_X1 port map( A1 => n15384, A2 => n15383, A3 => n15382, A4 => 
                           n15381, ZN => n15385);
   U13579 : NOR3_X1 port map( A1 => n15387, A2 => n15386, A3 => n15385, ZN => 
                           n15393);
   U13580 : AOI22_X1 port map( A1 => REGISTERS_5_55_port, A2 => n16518, B1 => 
                           REGISTERS_4_55_port, B2 => n16543, ZN => n15391);
   U13581 : AOI22_X1 port map( A1 => REGISTERS_7_55_port, A2 => n16594, B1 => 
                           REGISTERS_6_55_port, B2 => n16546, ZN => n15390);
   U13582 : AOI22_X1 port map( A1 => REGISTERS_0_55_port, A2 => n16597, B1 => 
                           REGISTERS_2_55_port, B2 => n16596, ZN => n15389);
   U13583 : AOI22_X1 port map( A1 => REGISTERS_3_55_port, A2 => n16453, B1 => 
                           REGISTERS_1_55_port, B2 => n16430, ZN => n15388);
   U13584 : AND4_X1 port map( A1 => n15391, A2 => n15390, A3 => n15389, A4 => 
                           n15388, ZN => n15392);
   U13585 : OAI222_X1 port map( A1 => n16605, A2 => n15393, B1 => n16553, B2 =>
                           n15392, C1 => n16026, C2 => n8433, ZN => n8578);
   U13586 : AOI22_X1 port map( A1 => REGISTERS_31_54_port, A2 => n16583, B1 => 
                           REGISTERS_23_54_port, B2 => n16572, ZN => n15397);
   U13587 : AOI22_X1 port map( A1 => REGISTERS_19_54_port, A2 => n16569, B1 => 
                           REGISTERS_20_54_port, B2 => n16581, ZN => n15396);
   U13588 : AOI22_X1 port map( A1 => REGISTERS_24_54_port, A2 => n16559, B1 => 
                           REGISTERS_30_54_port, B2 => n16555, ZN => n15395);
   U13589 : AOI22_X1 port map( A1 => REGISTERS_18_54_port, A2 => n16584, B1 => 
                           REGISTERS_22_54_port, B2 => n16556, ZN => n15394);
   U13590 : NAND4_X1 port map( A1 => n15397, A2 => n15396, A3 => n15395, A4 => 
                           n15394, ZN => n15408);
   U13591 : AOI22_X1 port map( A1 => REGISTERS_10_54_port, A2 => n16560, B1 => 
                           REGISTERS_29_54_port, B2 => n16574, ZN => n15401);
   U13592 : AOI22_X1 port map( A1 => REGISTERS_9_54_port, A2 => n16437, B1 => 
                           REGISTERS_21_54_port, B2 => n16568, ZN => n15400);
   U13593 : AOI22_X1 port map( A1 => REGISTERS_25_54_port, A2 => n16557, B1 => 
                           REGISTERS_27_54_port, B2 => n16573, ZN => n15399);
   U13594 : AOI22_X1 port map( A1 => REGISTERS_8_54_port, A2 => n16567, B1 => 
                           REGISTERS_15_54_port, B2 => n16558, ZN => n15398);
   U13595 : NAND4_X1 port map( A1 => n15401, A2 => n15400, A3 => n15399, A4 => 
                           n15398, ZN => n15407);
   U13596 : AOI22_X1 port map( A1 => REGISTERS_12_54_port, A2 => n16580, B1 => 
                           REGISTERS_13_54_port, B2 => n16562, ZN => n15405);
   U13597 : AOI22_X1 port map( A1 => REGISTERS_16_54_port, A2 => n16561, B1 => 
                           REGISTERS_26_54_port, B2 => n16582, ZN => n15404);
   U13598 : AOI22_X1 port map( A1 => REGISTERS_17_54_port, A2 => n16579, B1 => 
                           REGISTERS_11_54_port, B2 => n16414, ZN => n15403);
   U13599 : AOI22_X1 port map( A1 => REGISTERS_28_54_port, A2 => n16570, B1 => 
                           REGISTERS_14_54_port, B2 => n16571, ZN => n15402);
   U13600 : NAND4_X1 port map( A1 => n15405, A2 => n15404, A3 => n15403, A4 => 
                           n15402, ZN => n15406);
   U13601 : NOR3_X1 port map( A1 => n15408, A2 => n15407, A3 => n15406, ZN => 
                           n15414);
   U13602 : AOI22_X1 port map( A1 => REGISTERS_2_54_port, A2 => n16545, B1 => 
                           REGISTERS_4_54_port, B2 => n16543, ZN => n15412);
   U13603 : AOI22_X1 port map( A1 => REGISTERS_1_54_port, A2 => n16544, B1 => 
                           REGISTERS_6_54_port, B2 => n16546, ZN => n15411);
   U13604 : AOI22_X1 port map( A1 => REGISTERS_5_54_port, A2 => n16542, B1 => 
                           REGISTERS_0_54_port, B2 => n16597, ZN => n15410);
   U13605 : AOI22_X1 port map( A1 => REGISTERS_3_54_port, A2 => n16453, B1 => 
                           REGISTERS_7_54_port, B2 => n16594, ZN => n15409);
   U13606 : AND4_X1 port map( A1 => n15412, A2 => n15411, A3 => n15410, A4 => 
                           n15409, ZN => n15413);
   U13607 : OAI222_X1 port map( A1 => n16605, A2 => n15414, B1 => n16603, B2 =>
                           n15413, C1 => n16026, C2 => n8432, ZN => n8579);
   U13608 : AOI22_X1 port map( A1 => REGISTERS_21_53_port, A2 => n16568, B1 => 
                           REGISTERS_10_53_port, B2 => n16560, ZN => n15418);
   U13609 : AOI22_X1 port map( A1 => REGISTERS_8_53_port, A2 => n16567, B1 => 
                           REGISTERS_30_53_port, B2 => n16555, ZN => n15417);
   U13610 : AOI22_X1 port map( A1 => REGISTERS_18_53_port, A2 => n16584, B1 => 
                           REGISTERS_31_53_port, B2 => n16583, ZN => n15416);
   U13611 : AOI22_X1 port map( A1 => REGISTERS_9_53_port, A2 => n16029, B1 => 
                           REGISTERS_28_53_port, B2 => n16570, ZN => n15415);
   U13612 : NAND4_X1 port map( A1 => n15418, A2 => n15417, A3 => n15416, A4 => 
                           n15415, ZN => n15429);
   U13613 : AOI22_X1 port map( A1 => REGISTERS_20_53_port, A2 => n16581, B1 => 
                           REGISTERS_29_53_port, B2 => n16574, ZN => n15422);
   U13614 : AOI22_X1 port map( A1 => REGISTERS_14_53_port, A2 => n16571, B1 => 
                           REGISTERS_17_53_port, B2 => n16579, ZN => n15421);
   U13615 : AOI22_X1 port map( A1 => REGISTERS_23_53_port, A2 => n16572, B1 => 
                           REGISTERS_27_53_port, B2 => n16573, ZN => n15420);
   U13616 : AOI22_X1 port map( A1 => REGISTERS_13_53_port, A2 => n16562, B1 => 
                           REGISTERS_12_53_port, B2 => n16580, ZN => n15419);
   U13617 : NAND4_X1 port map( A1 => n15422, A2 => n15421, A3 => n15420, A4 => 
                           n15419, ZN => n15428);
   U13618 : AOI22_X1 port map( A1 => REGISTERS_26_53_port, A2 => n16582, B1 => 
                           REGISTERS_25_53_port, B2 => n16557, ZN => n15426);
   U13619 : AOI22_X1 port map( A1 => REGISTERS_22_53_port, A2 => n16556, B1 => 
                           REGISTERS_19_53_port, B2 => n16569, ZN => n15425);
   U13620 : AOI22_X1 port map( A1 => REGISTERS_16_53_port, A2 => n16561, B1 => 
                           REGISTERS_24_53_port, B2 => n16559, ZN => n15424);
   U13621 : AOI22_X1 port map( A1 => REGISTERS_15_53_port, A2 => n16558, B1 => 
                           REGISTERS_11_53_port, B2 => n16414, ZN => n15423);
   U13622 : NAND4_X1 port map( A1 => n15426, A2 => n15425, A3 => n15424, A4 => 
                           n15423, ZN => n15427);
   U13623 : NOR3_X1 port map( A1 => n15429, A2 => n15428, A3 => n15427, ZN => 
                           n15435);
   U13624 : AOI22_X1 port map( A1 => REGISTERS_0_53_port, A2 => n16597, B1 => 
                           REGISTERS_1_53_port, B2 => n16430, ZN => n15433);
   U13625 : AOI22_X1 port map( A1 => REGISTERS_2_53_port, A2 => n16596, B1 => 
                           REGISTERS_3_53_port, B2 => n16593, ZN => n15432);
   U13626 : AOI22_X1 port map( A1 => REGISTERS_6_53_port, A2 => n16546, B1 => 
                           REGISTERS_5_53_port, B2 => n16542, ZN => n15431);
   U13627 : AOI22_X1 port map( A1 => REGISTERS_4_53_port, A2 => n16595, B1 => 
                           REGISTERS_7_53_port, B2 => n16454, ZN => n15430);
   U13628 : AND4_X1 port map( A1 => n15433, A2 => n15432, A3 => n15431, A4 => 
                           n15430, ZN => n15434);
   U13629 : OAI222_X1 port map( A1 => n15796, A2 => n15435, B1 => n16553, B2 =>
                           n15434, C1 => n16049, C2 => n8431, ZN => n8580);
   U13630 : AOI22_X1 port map( A1 => REGISTERS_12_52_port, A2 => n16580, B1 => 
                           REGISTERS_20_52_port, B2 => n16581, ZN => n15439);
   U13631 : AOI22_X1 port map( A1 => REGISTERS_14_52_port, A2 => n16571, B1 => 
                           REGISTERS_27_52_port, B2 => n16573, ZN => n15438);
   U13632 : AOI22_X1 port map( A1 => REGISTERS_17_52_port, A2 => n16579, B1 => 
                           REGISTERS_21_52_port, B2 => n16568, ZN => n15437);
   U13633 : AOI22_X1 port map( A1 => REGISTERS_16_52_port, A2 => n16561, B1 => 
                           REGISTERS_28_52_port, B2 => n16570, ZN => n15436);
   U13634 : NAND4_X1 port map( A1 => n15439, A2 => n15438, A3 => n15437, A4 => 
                           n15436, ZN => n15450);
   U13635 : AOI22_X1 port map( A1 => REGISTERS_22_52_port, A2 => n16556, B1 => 
                           REGISTERS_30_52_port, B2 => n16555, ZN => n15443);
   U13636 : AOI22_X1 port map( A1 => REGISTERS_26_52_port, A2 => n16582, B1 => 
                           REGISTERS_25_52_port, B2 => n16557, ZN => n15442);
   U13637 : AOI22_X1 port map( A1 => REGISTERS_15_52_port, A2 => n16558, B1 => 
                           REGISTERS_8_52_port, B2 => n16567, ZN => n15441);
   U13638 : AOI22_X1 port map( A1 => REGISTERS_13_52_port, A2 => n16562, B1 => 
                           REGISTERS_19_52_port, B2 => n16569, ZN => n15440);
   U13639 : NAND4_X1 port map( A1 => n15443, A2 => n15442, A3 => n15441, A4 => 
                           n15440, ZN => n15449);
   U13640 : AOI22_X1 port map( A1 => REGISTERS_9_52_port, A2 => n16437, B1 => 
                           REGISTERS_31_52_port, B2 => n16583, ZN => n15447);
   U13641 : AOI22_X1 port map( A1 => REGISTERS_24_52_port, A2 => n16559, B1 => 
                           REGISTERS_29_52_port, B2 => n16574, ZN => n15446);
   U13642 : AOI22_X1 port map( A1 => REGISTERS_18_52_port, A2 => n16584, B1 => 
                           REGISTERS_11_52_port, B2 => n15782, ZN => n15445);
   U13643 : AOI22_X1 port map( A1 => REGISTERS_23_52_port, A2 => n16572, B1 => 
                           REGISTERS_10_52_port, B2 => n16560, ZN => n15444);
   U13644 : NAND4_X1 port map( A1 => n15447, A2 => n15446, A3 => n15445, A4 => 
                           n15444, ZN => n15448);
   U13645 : NOR3_X1 port map( A1 => n15450, A2 => n15449, A3 => n15448, ZN => 
                           n15456);
   U13646 : AOI22_X1 port map( A1 => REGISTERS_5_52_port, A2 => n16518, B1 => 
                           REGISTERS_1_52_port, B2 => n16544, ZN => n15454);
   U13647 : AOI22_X1 port map( A1 => REGISTERS_7_52_port, A2 => n16454, B1 => 
                           REGISTERS_6_52_port, B2 => n16592, ZN => n15453);
   U13648 : AOI22_X1 port map( A1 => REGISTERS_3_52_port, A2 => n16453, B1 => 
                           REGISTERS_2_52_port, B2 => n16545, ZN => n15452);
   U13649 : AOI22_X1 port map( A1 => REGISTERS_0_52_port, A2 => n16597, B1 => 
                           REGISTERS_4_52_port, B2 => n16543, ZN => n15451);
   U13650 : AND4_X1 port map( A1 => n15454, A2 => n15453, A3 => n15452, A4 => 
                           n15451, ZN => n15455);
   U13651 : OAI222_X1 port map( A1 => n16605, A2 => n15456, B1 => n16603, B2 =>
                           n15455, C1 => n16026, C2 => n8430, ZN => n8581);
   U13652 : AOI22_X1 port map( A1 => REGISTERS_30_51_port, A2 => n16555, B1 => 
                           REGISTERS_13_51_port, B2 => n16562, ZN => n15460);
   U13653 : AOI22_X1 port map( A1 => REGISTERS_21_51_port, A2 => n16568, B1 => 
                           REGISTERS_22_51_port, B2 => n16556, ZN => n15459);
   U13654 : AOI22_X1 port map( A1 => REGISTERS_14_51_port, A2 => n16571, B1 => 
                           REGISTERS_12_51_port, B2 => n16580, ZN => n15458);
   U13655 : AOI22_X1 port map( A1 => REGISTERS_28_51_port, A2 => n16570, B1 => 
                           REGISTERS_25_51_port, B2 => n16557, ZN => n15457);
   U13656 : NAND4_X1 port map( A1 => n15460, A2 => n15459, A3 => n15458, A4 => 
                           n15457, ZN => n15471);
   U13657 : AOI22_X1 port map( A1 => REGISTERS_26_51_port, A2 => n16582, B1 => 
                           REGISTERS_31_51_port, B2 => n16583, ZN => n15464);
   U13658 : AOI22_X1 port map( A1 => REGISTERS_18_51_port, A2 => n16584, B1 => 
                           REGISTERS_29_51_port, B2 => n16574, ZN => n15463);
   U13659 : AOI22_X1 port map( A1 => REGISTERS_19_51_port, A2 => n16569, B1 => 
                           REGISTERS_10_51_port, B2 => n16560, ZN => n15462);
   U13660 : AOI22_X1 port map( A1 => REGISTERS_24_51_port, A2 => n16559, B1 => 
                           REGISTERS_20_51_port, B2 => n16581, ZN => n15461);
   U13661 : NAND4_X1 port map( A1 => n15464, A2 => n15463, A3 => n15462, A4 => 
                           n15461, ZN => n15470);
   U13662 : AOI22_X1 port map( A1 => REGISTERS_23_51_port, A2 => n16572, B1 => 
                           REGISTERS_16_51_port, B2 => n16561, ZN => n15468);
   U13663 : AOI22_X1 port map( A1 => REGISTERS_11_51_port, A2 => n16414, B1 => 
                           REGISTERS_9_51_port, B2 => n16029, ZN => n15467);
   U13664 : AOI22_X1 port map( A1 => REGISTERS_8_51_port, A2 => n16567, B1 => 
                           REGISTERS_27_51_port, B2 => n16573, ZN => n15466);
   U13665 : AOI22_X1 port map( A1 => REGISTERS_17_51_port, A2 => n16579, B1 => 
                           REGISTERS_15_51_port, B2 => n16558, ZN => n15465);
   U13666 : NAND4_X1 port map( A1 => n15468, A2 => n15467, A3 => n15466, A4 => 
                           n15465, ZN => n15469);
   U13667 : NOR3_X1 port map( A1 => n15471, A2 => n15470, A3 => n15469, ZN => 
                           n15477);
   U13668 : AOI22_X1 port map( A1 => REGISTERS_6_51_port, A2 => n16592, B1 => 
                           REGISTERS_0_51_port, B2 => n16547, ZN => n15475);
   U13669 : AOI22_X1 port map( A1 => REGISTERS_3_51_port, A2 => n16453, B1 => 
                           REGISTERS_5_51_port, B2 => n16518, ZN => n15474);
   U13670 : AOI22_X1 port map( A1 => REGISTERS_2_51_port, A2 => n16545, B1 => 
                           REGISTERS_1_51_port, B2 => n16430, ZN => n15473);
   U13671 : AOI22_X1 port map( A1 => REGISTERS_7_51_port, A2 => n16594, B1 => 
                           REGISTERS_4_51_port, B2 => n16595, ZN => n15472);
   U13672 : AND4_X1 port map( A1 => n15475, A2 => n15474, A3 => n15473, A4 => 
                           n15472, ZN => n15476);
   U13673 : OAI222_X1 port map( A1 => n15796, A2 => n15477, B1 => n16553, B2 =>
                           n15476, C1 => n16026, C2 => n8429, ZN => n8582);
   U13674 : AOI22_X1 port map( A1 => REGISTERS_24_50_port, A2 => n16559, B1 => 
                           REGISTERS_29_50_port, B2 => n16574, ZN => n15481);
   U13675 : AOI22_X1 port map( A1 => REGISTERS_27_50_port, A2 => n16573, B1 => 
                           REGISTERS_16_50_port, B2 => n16561, ZN => n15480);
   U13676 : AOI22_X1 port map( A1 => REGISTERS_31_50_port, A2 => n16583, B1 => 
                           REGISTERS_23_50_port, B2 => n16572, ZN => n15479);
   U13677 : AOI22_X1 port map( A1 => REGISTERS_28_50_port, A2 => n16570, B1 => 
                           REGISTERS_11_50_port, B2 => n15782, ZN => n15478);
   U13678 : NAND4_X1 port map( A1 => n15481, A2 => n15480, A3 => n15479, A4 => 
                           n15478, ZN => n15492);
   U13679 : AOI22_X1 port map( A1 => REGISTERS_25_50_port, A2 => n16557, B1 => 
                           REGISTERS_22_50_port, B2 => n16556, ZN => n15485);
   U13680 : AOI22_X1 port map( A1 => REGISTERS_17_50_port, A2 => n16579, B1 => 
                           REGISTERS_19_50_port, B2 => n16569, ZN => n15484);
   U13681 : AOI22_X1 port map( A1 => REGISTERS_26_50_port, A2 => n16582, B1 => 
                           REGISTERS_21_50_port, B2 => n16568, ZN => n15483);
   U13682 : AOI22_X1 port map( A1 => REGISTERS_8_50_port, A2 => n16567, B1 => 
                           REGISTERS_12_50_port, B2 => n16580, ZN => n15482);
   U13683 : NAND4_X1 port map( A1 => n15485, A2 => n15484, A3 => n15483, A4 => 
                           n15482, ZN => n15491);
   U13684 : AOI22_X1 port map( A1 => REGISTERS_30_50_port, A2 => n16555, B1 => 
                           REGISTERS_15_50_port, B2 => n16558, ZN => n15489);
   U13685 : AOI22_X1 port map( A1 => REGISTERS_14_50_port, A2 => n16571, B1 => 
                           REGISTERS_20_50_port, B2 => n16581, ZN => n15488);
   U13686 : AOI22_X1 port map( A1 => REGISTERS_10_50_port, A2 => n16560, B1 => 
                           REGISTERS_18_50_port, B2 => n16584, ZN => n15487);
   U13687 : AOI22_X1 port map( A1 => REGISTERS_13_50_port, A2 => n16562, B1 => 
                           REGISTERS_9_50_port, B2 => n16029, ZN => n15486);
   U13688 : NAND4_X1 port map( A1 => n15489, A2 => n15488, A3 => n15487, A4 => 
                           n15486, ZN => n15490);
   U13689 : NOR3_X1 port map( A1 => n15492, A2 => n15491, A3 => n15490, ZN => 
                           n15498);
   U13690 : AOI22_X1 port map( A1 => REGISTERS_5_50_port, A2 => n16542, B1 => 
                           REGISTERS_6_50_port, B2 => n16592, ZN => n15496);
   U13691 : AOI22_X1 port map( A1 => REGISTERS_1_50_port, A2 => n16544, B1 => 
                           REGISTERS_7_50_port, B2 => n16594, ZN => n15495);
   U13692 : AOI22_X1 port map( A1 => REGISTERS_3_50_port, A2 => n16453, B1 => 
                           REGISTERS_4_50_port, B2 => n16543, ZN => n15494);
   U13693 : AOI22_X1 port map( A1 => REGISTERS_2_50_port, A2 => n16596, B1 => 
                           REGISTERS_0_50_port, B2 => n16547, ZN => n15493);
   U13694 : AND4_X1 port map( A1 => n15496, A2 => n15495, A3 => n15494, A4 => 
                           n15493, ZN => n15497);
   U13695 : OAI222_X1 port map( A1 => n15796, A2 => n15498, B1 => n16553, B2 =>
                           n15497, C1 => n16026, C2 => n8428, ZN => n8583);
   U13696 : AOI22_X1 port map( A1 => REGISTERS_8_49_port, A2 => n16567, B1 => 
                           REGISTERS_11_49_port, B2 => n15782, ZN => n15502);
   U13697 : AOI22_X1 port map( A1 => REGISTERS_17_49_port, A2 => n16579, B1 => 
                           REGISTERS_15_49_port, B2 => n16558, ZN => n15501);
   U13698 : AOI22_X1 port map( A1 => REGISTERS_9_49_port, A2 => n16525, B1 => 
                           REGISTERS_10_49_port, B2 => n16560, ZN => n15500);
   U13699 : AOI22_X1 port map( A1 => REGISTERS_28_49_port, A2 => n16570, B1 => 
                           REGISTERS_27_49_port, B2 => n16573, ZN => n15499);
   U13700 : NAND4_X1 port map( A1 => n15502, A2 => n15501, A3 => n15500, A4 => 
                           n15499, ZN => n15513);
   U13701 : AOI22_X1 port map( A1 => REGISTERS_13_49_port, A2 => n16562, B1 => 
                           REGISTERS_19_49_port, B2 => n16569, ZN => n15506);
   U13702 : AOI22_X1 port map( A1 => REGISTERS_25_49_port, A2 => n16557, B1 => 
                           REGISTERS_22_49_port, B2 => n16556, ZN => n15505);
   U13703 : AOI22_X1 port map( A1 => REGISTERS_23_49_port, A2 => n16572, B1 => 
                           REGISTERS_20_49_port, B2 => n16581, ZN => n15504);
   U13704 : AOI22_X1 port map( A1 => REGISTERS_21_49_port, A2 => n16568, B1 => 
                           REGISTERS_18_49_port, B2 => n16584, ZN => n15503);
   U13705 : NAND4_X1 port map( A1 => n15506, A2 => n15505, A3 => n15504, A4 => 
                           n15503, ZN => n15512);
   U13706 : AOI22_X1 port map( A1 => REGISTERS_24_49_port, A2 => n16559, B1 => 
                           REGISTERS_14_49_port, B2 => n16571, ZN => n15510);
   U13707 : AOI22_X1 port map( A1 => REGISTERS_31_49_port, A2 => n16583, B1 => 
                           REGISTERS_29_49_port, B2 => n16574, ZN => n15509);
   U13708 : AOI22_X1 port map( A1 => REGISTERS_26_49_port, A2 => n16582, B1 => 
                           REGISTERS_16_49_port, B2 => n16561, ZN => n15508);
   U13709 : AOI22_X1 port map( A1 => REGISTERS_30_49_port, A2 => n16555, B1 => 
                           REGISTERS_12_49_port, B2 => n16580, ZN => n15507);
   U13710 : NAND4_X1 port map( A1 => n15510, A2 => n15509, A3 => n15508, A4 => 
                           n15507, ZN => n15511);
   U13711 : NOR3_X1 port map( A1 => n15513, A2 => n15512, A3 => n15511, ZN => 
                           n15519);
   U13712 : AOI22_X1 port map( A1 => REGISTERS_7_49_port, A2 => n16594, B1 => 
                           REGISTERS_5_49_port, B2 => n16542, ZN => n15517);
   U13713 : AOI22_X1 port map( A1 => REGISTERS_3_49_port, A2 => n16453, B1 => 
                           REGISTERS_4_49_port, B2 => n16595, ZN => n15516);
   U13714 : AOI22_X1 port map( A1 => REGISTERS_6_49_port, A2 => n16592, B1 => 
                           REGISTERS_2_49_port, B2 => n16596, ZN => n15515);
   U13715 : AOI22_X1 port map( A1 => REGISTERS_1_49_port, A2 => n16544, B1 => 
                           REGISTERS_0_49_port, B2 => n16547, ZN => n15514);
   U13716 : OAI222_X1 port map( A1 => n16605, A2 => n15519, B1 => n16553, B2 =>
                           n15518, C1 => n16049, C2 => n8427, ZN => n8584);
   U13717 : AOI22_X1 port map( A1 => REGISTERS_23_48_port, A2 => n16572, B1 => 
                           REGISTERS_27_48_port, B2 => n16573, ZN => n15523);
   U13718 : AOI22_X1 port map( A1 => REGISTERS_10_48_port, A2 => n16560, B1 => 
                           REGISTERS_15_48_port, B2 => n16558, ZN => n15522);
   U13719 : AOI22_X1 port map( A1 => REGISTERS_25_48_port, A2 => n16557, B1 => 
                           REGISTERS_11_48_port, B2 => n15782, ZN => n15521);
   U13720 : AOI22_X1 port map( A1 => REGISTERS_20_48_port, A2 => n16581, B1 => 
                           REGISTERS_29_48_port, B2 => n16574, ZN => n15520);
   U13721 : NAND4_X1 port map( A1 => n15523, A2 => n15522, A3 => n15521, A4 => 
                           n15520, ZN => n15534);
   U13722 : AOI22_X1 port map( A1 => REGISTERS_17_48_port, A2 => n16579, B1 => 
                           REGISTERS_18_48_port, B2 => n16584, ZN => n15527);
   U13723 : AOI22_X1 port map( A1 => REGISTERS_28_48_port, A2 => n16570, B1 => 
                           REGISTERS_21_48_port, B2 => n16568, ZN => n15526);
   U13724 : AOI22_X1 port map( A1 => REGISTERS_13_48_port, A2 => n16562, B1 => 
                           REGISTERS_19_48_port, B2 => n16569, ZN => n15525);
   U13725 : AOI22_X1 port map( A1 => REGISTERS_8_48_port, A2 => n16567, B1 => 
                           REGISTERS_22_48_port, B2 => n16556, ZN => n15524);
   U13726 : NAND4_X1 port map( A1 => n15527, A2 => n15526, A3 => n15525, A4 => 
                           n15524, ZN => n15533);
   U13727 : AOI22_X1 port map( A1 => REGISTERS_31_48_port, A2 => n16583, B1 => 
                           REGISTERS_26_48_port, B2 => n16582, ZN => n15531);
   U13728 : AOI22_X1 port map( A1 => REGISTERS_12_48_port, A2 => n16580, B1 => 
                           REGISTERS_9_48_port, B2 => n16029, ZN => n15530);
   U13729 : AOI22_X1 port map( A1 => REGISTERS_24_48_port, A2 => n16559, B1 => 
                           REGISTERS_30_48_port, B2 => n16555, ZN => n15529);
   U13730 : AOI22_X1 port map( A1 => REGISTERS_14_48_port, A2 => n16571, B1 => 
                           REGISTERS_16_48_port, B2 => n16561, ZN => n15528);
   U13731 : NAND4_X1 port map( A1 => n15531, A2 => n15530, A3 => n15529, A4 => 
                           n15528, ZN => n15532);
   U13732 : NOR3_X1 port map( A1 => n15534, A2 => n15533, A3 => n15532, ZN => 
                           n15540);
   U13733 : AOI22_X1 port map( A1 => REGISTERS_1_48_port, A2 => n16430, B1 => 
                           REGISTERS_7_48_port, B2 => n16594, ZN => n15538);
   U13734 : AOI22_X1 port map( A1 => REGISTERS_2_48_port, A2 => n16545, B1 => 
                           REGISTERS_4_48_port, B2 => n16543, ZN => n15537);
   U13735 : AOI22_X1 port map( A1 => REGISTERS_6_48_port, A2 => n16546, B1 => 
                           REGISTERS_5_48_port, B2 => n16542, ZN => n15536);
   U13736 : AOI22_X1 port map( A1 => REGISTERS_0_48_port, A2 => n16597, B1 => 
                           REGISTERS_3_48_port, B2 => n16453, ZN => n15535);
   U13737 : AND4_X1 port map( A1 => n15538, A2 => n15537, A3 => n15536, A4 => 
                           n15535, ZN => n15539);
   U13738 : OAI222_X1 port map( A1 => n16605, A2 => n15540, B1 => n16553, B2 =>
                           n15539, C1 => n16026, C2 => n8426, ZN => n8585);
   U13739 : AOI22_X1 port map( A1 => REGISTERS_23_47_port, A2 => n16572, B1 => 
                           REGISTERS_10_47_port, B2 => n16560, ZN => n15544);
   U13740 : AOI22_X1 port map( A1 => REGISTERS_20_47_port, A2 => n16581, B1 => 
                           REGISTERS_11_47_port, B2 => n15782, ZN => n15543);
   U13741 : AOI22_X1 port map( A1 => REGISTERS_8_47_port, A2 => n16567, B1 => 
                           REGISTERS_28_47_port, B2 => n16570, ZN => n15542);
   U13742 : AOI22_X1 port map( A1 => REGISTERS_17_47_port, A2 => n16579, B1 => 
                           REGISTERS_31_47_port, B2 => n16583, ZN => n15541);
   U13743 : NAND4_X1 port map( A1 => n15544, A2 => n15543, A3 => n15542, A4 => 
                           n15541, ZN => n15555);
   U13744 : AOI22_X1 port map( A1 => REGISTERS_14_47_port, A2 => n16571, B1 => 
                           REGISTERS_15_47_port, B2 => n16558, ZN => n15548);
   U13745 : AOI22_X1 port map( A1 => REGISTERS_18_47_port, A2 => n16584, B1 => 
                           REGISTERS_16_47_port, B2 => n16561, ZN => n15547);
   U13746 : AOI22_X1 port map( A1 => REGISTERS_27_47_port, A2 => n16573, B1 => 
                           REGISTERS_25_47_port, B2 => n16557, ZN => n15546);
   U13747 : AOI22_X1 port map( A1 => REGISTERS_13_47_port, A2 => n16562, B1 => 
                           REGISTERS_29_47_port, B2 => n16574, ZN => n15545);
   U13748 : NAND4_X1 port map( A1 => n15548, A2 => n15547, A3 => n15546, A4 => 
                           n15545, ZN => n15554);
   U13749 : AOI22_X1 port map( A1 => REGISTERS_21_47_port, A2 => n16568, B1 => 
                           REGISTERS_30_47_port, B2 => n16555, ZN => n15552);
   U13750 : AOI22_X1 port map( A1 => REGISTERS_26_47_port, A2 => n16582, B1 => 
                           REGISTERS_24_47_port, B2 => n16559, ZN => n15551);
   U13751 : AOI22_X1 port map( A1 => REGISTERS_22_47_port, A2 => n16556, B1 => 
                           REGISTERS_9_47_port, B2 => n16029, ZN => n15550);
   U13752 : AOI22_X1 port map( A1 => REGISTERS_19_47_port, A2 => n16569, B1 => 
                           REGISTERS_12_47_port, B2 => n16580, ZN => n15549);
   U13753 : NAND4_X1 port map( A1 => n15552, A2 => n15551, A3 => n15550, A4 => 
                           n15549, ZN => n15553);
   U13754 : NOR3_X1 port map( A1 => n15555, A2 => n15554, A3 => n15553, ZN => 
                           n15562);
   U13755 : AOI22_X1 port map( A1 => REGISTERS_5_47_port, A2 => n16518, B1 => 
                           REGISTERS_6_47_port, B2 => n16592, ZN => n15560);
   U13756 : AOI22_X1 port map( A1 => REGISTERS_0_47_port, A2 => n16547, B1 => 
                           REGISTERS_1_47_port, B2 => n16430, ZN => n15559);
   U13757 : AOI22_X1 port map( A1 => REGISTERS_4_47_port, A2 => n16543, B1 => 
                           REGISTERS_7_47_port, B2 => n16594, ZN => n15558);
   U13758 : AOI22_X1 port map( A1 => REGISTERS_3_47_port, A2 => n16453, B1 => 
                           REGISTERS_2_47_port, B2 => n16545, ZN => n15557);
   U13759 : AND4_X1 port map( A1 => n15560, A2 => n15559, A3 => n15558, A4 => 
                           n15557, ZN => n15561);
   U13760 : OAI222_X1 port map( A1 => n15796, A2 => n15562, B1 => n16553, B2 =>
                           n15561, C1 => n16026, C2 => n8425, ZN => n8586);
   U13761 : AOI22_X1 port map( A1 => REGISTERS_8_46_port, A2 => n16567, B1 => 
                           REGISTERS_14_46_port, B2 => n16571, ZN => n15566);
   U13762 : AOI22_X1 port map( A1 => REGISTERS_27_46_port, A2 => n16573, B1 => 
                           REGISTERS_26_46_port, B2 => n16582, ZN => n15565);
   U13763 : AOI22_X1 port map( A1 => REGISTERS_18_46_port, A2 => n16584, B1 => 
                           REGISTERS_16_46_port, B2 => n16561, ZN => n15564);
   U13764 : AOI22_X1 port map( A1 => REGISTERS_15_46_port, A2 => n16558, B1 => 
                           REGISTERS_19_46_port, B2 => n16569, ZN => n15563);
   U13765 : NAND4_X1 port map( A1 => n15566, A2 => n15565, A3 => n15564, A4 => 
                           n15563, ZN => n15577);
   U13766 : AOI22_X1 port map( A1 => REGISTERS_17_46_port, A2 => n16579, B1 => 
                           REGISTERS_20_46_port, B2 => n16581, ZN => n15570);
   U13767 : AOI22_X1 port map( A1 => REGISTERS_23_46_port, A2 => n16572, B1 => 
                           REGISTERS_30_46_port, B2 => n16555, ZN => n15569);
   U13768 : AOI22_X1 port map( A1 => REGISTERS_24_46_port, A2 => n16559, B1 => 
                           REGISTERS_11_46_port, B2 => n15782, ZN => n15568);
   U13769 : AOI22_X1 port map( A1 => REGISTERS_13_46_port, A2 => n16562, B1 => 
                           REGISTERS_10_46_port, B2 => n16560, ZN => n15567);
   U13770 : NAND4_X1 port map( A1 => n15570, A2 => n15569, A3 => n15568, A4 => 
                           n15567, ZN => n15576);
   U13771 : AOI22_X1 port map( A1 => REGISTERS_12_46_port, A2 => n16580, B1 => 
                           REGISTERS_31_46_port, B2 => n16583, ZN => n15574);
   U13772 : AOI22_X1 port map( A1 => REGISTERS_9_46_port, A2 => n16525, B1 => 
                           REGISTERS_29_46_port, B2 => n16574, ZN => n15573);
   U13773 : AOI22_X1 port map( A1 => REGISTERS_25_46_port, A2 => n16557, B1 => 
                           REGISTERS_28_46_port, B2 => n16570, ZN => n15572);
   U13774 : AOI22_X1 port map( A1 => REGISTERS_21_46_port, A2 => n16568, B1 => 
                           REGISTERS_22_46_port, B2 => n16556, ZN => n15571);
   U13775 : NAND4_X1 port map( A1 => n15574, A2 => n15573, A3 => n15572, A4 => 
                           n15571, ZN => n15575);
   U13776 : NOR3_X1 port map( A1 => n15577, A2 => n15576, A3 => n15575, ZN => 
                           n15583);
   U13777 : AOI22_X1 port map( A1 => REGISTERS_3_46_port, A2 => n15746, B1 => 
                           REGISTERS_7_46_port, B2 => n16594, ZN => n15581);
   U13778 : AOI22_X1 port map( A1 => REGISTERS_2_46_port, A2 => n16545, B1 => 
                           REGISTERS_4_46_port, B2 => n16595, ZN => n15580);
   U13779 : AOI22_X1 port map( A1 => REGISTERS_5_46_port, A2 => n16542, B1 => 
                           REGISTERS_0_46_port, B2 => n16547, ZN => n15579);
   U13780 : AOI22_X1 port map( A1 => REGISTERS_6_46_port, A2 => n16592, B1 => 
                           REGISTERS_1_46_port, B2 => n16544, ZN => n15578);
   U13781 : AND4_X1 port map( A1 => n15581, A2 => n15580, A3 => n15579, A4 => 
                           n15578, ZN => n15582);
   U13782 : OAI222_X1 port map( A1 => n15796, A2 => n15583, B1 => n16553, B2 =>
                           n15582, C1 => n16026, C2 => n8424, ZN => n8587);
   U13783 : AOI22_X1 port map( A1 => REGISTERS_16_45_port, A2 => n16561, B1 => 
                           REGISTERS_20_45_port, B2 => n16581, ZN => n15587);
   U13784 : AOI22_X1 port map( A1 => REGISTERS_18_45_port, A2 => n16584, B1 => 
                           REGISTERS_28_45_port, B2 => n16570, ZN => n15586);
   U13785 : AOI22_X1 port map( A1 => REGISTERS_21_45_port, A2 => n16568, B1 => 
                           REGISTERS_31_45_port, B2 => n16583, ZN => n15585);
   U13786 : AOI22_X1 port map( A1 => REGISTERS_17_45_port, A2 => n16579, B1 => 
                           REGISTERS_14_45_port, B2 => n16571, ZN => n15584);
   U13787 : NAND4_X1 port map( A1 => n15587, A2 => n15586, A3 => n15585, A4 => 
                           n15584, ZN => n15598);
   U13788 : AOI22_X1 port map( A1 => REGISTERS_12_45_port, A2 => n16580, B1 => 
                           REGISTERS_11_45_port, B2 => n15782, ZN => n15591);
   U13789 : AOI22_X1 port map( A1 => REGISTERS_25_45_port, A2 => n16557, B1 => 
                           REGISTERS_15_45_port, B2 => n16558, ZN => n15590);
   U13790 : AOI22_X1 port map( A1 => REGISTERS_9_45_port, A2 => n16029, B1 => 
                           REGISTERS_24_45_port, B2 => n16559, ZN => n15589);
   U13791 : AOI22_X1 port map( A1 => REGISTERS_29_45_port, A2 => n16574, B1 => 
                           REGISTERS_19_45_port, B2 => n16569, ZN => n15588);
   U13792 : NAND4_X1 port map( A1 => n15591, A2 => n15590, A3 => n15589, A4 => 
                           n15588, ZN => n15597);
   U13793 : AOI22_X1 port map( A1 => REGISTERS_22_45_port, A2 => n16556, B1 => 
                           REGISTERS_27_45_port, B2 => n16573, ZN => n15595);
   U13794 : AOI22_X1 port map( A1 => REGISTERS_10_45_port, A2 => n16560, B1 => 
                           REGISTERS_30_45_port, B2 => n16555, ZN => n15594);
   U13795 : AOI22_X1 port map( A1 => REGISTERS_8_45_port, A2 => n16567, B1 => 
                           REGISTERS_26_45_port, B2 => n16582, ZN => n15593);
   U13796 : AOI22_X1 port map( A1 => REGISTERS_13_45_port, A2 => n16562, B1 => 
                           REGISTERS_23_45_port, B2 => n16572, ZN => n15592);
   U13797 : NAND4_X1 port map( A1 => n15595, A2 => n15594, A3 => n15593, A4 => 
                           n15592, ZN => n15596);
   U13798 : NOR3_X1 port map( A1 => n15598, A2 => n15597, A3 => n15596, ZN => 
                           n15604);
   U13799 : AOI22_X1 port map( A1 => REGISTERS_1_45_port, A2 => n16544, B1 => 
                           REGISTERS_7_45_port, B2 => n16594, ZN => n15602);
   U13800 : AOI22_X1 port map( A1 => REGISTERS_0_45_port, A2 => n16597, B1 => 
                           REGISTERS_4_45_port, B2 => n16595, ZN => n15601);
   U13801 : AOI22_X1 port map( A1 => REGISTERS_2_45_port, A2 => n16545, B1 => 
                           REGISTERS_6_45_port, B2 => n16546, ZN => n15600);
   U13802 : AOI22_X1 port map( A1 => REGISTERS_3_45_port, A2 => n15746, B1 => 
                           REGISTERS_5_45_port, B2 => n16518, ZN => n15599);
   U13803 : AND4_X1 port map( A1 => n15602, A2 => n15601, A3 => n15600, A4 => 
                           n15599, ZN => n15603);
   U13804 : OAI222_X1 port map( A1 => n15796, A2 => n15604, B1 => n16553, B2 =>
                           n15603, C1 => n16049, C2 => n8423, ZN => n8588);
   U13805 : AOI22_X1 port map( A1 => REGISTERS_19_44_port, A2 => n16569, B1 => 
                           REGISTERS_13_44_port, B2 => n16562, ZN => n15608);
   U13806 : AOI22_X1 port map( A1 => REGISTERS_17_44_port, A2 => n16579, B1 => 
                           REGISTERS_14_44_port, B2 => n16571, ZN => n15607);
   U13807 : AOI22_X1 port map( A1 => REGISTERS_8_44_port, A2 => n16567, B1 => 
                           REGISTERS_24_44_port, B2 => n16559, ZN => n15606);
   U13808 : AOI22_X1 port map( A1 => REGISTERS_20_44_port, A2 => n16581, B1 => 
                           REGISTERS_12_44_port, B2 => n16580, ZN => n15605);
   U13809 : NAND4_X1 port map( A1 => n15608, A2 => n15607, A3 => n15606, A4 => 
                           n15605, ZN => n15619);
   U13810 : AOI22_X1 port map( A1 => REGISTERS_25_44_port, A2 => n16557, B1 => 
                           REGISTERS_30_44_port, B2 => n16555, ZN => n15612);
   U13811 : AOI22_X1 port map( A1 => REGISTERS_21_44_port, A2 => n16568, B1 => 
                           REGISTERS_15_44_port, B2 => n16558, ZN => n15611);
   U13812 : AOI22_X1 port map( A1 => REGISTERS_27_44_port, A2 => n16573, B1 => 
                           REGISTERS_11_44_port, B2 => n15782, ZN => n15610);
   U13813 : AOI22_X1 port map( A1 => REGISTERS_18_44_port, A2 => n16584, B1 => 
                           REGISTERS_23_44_port, B2 => n16572, ZN => n15609);
   U13814 : NAND4_X1 port map( A1 => n15612, A2 => n15611, A3 => n15610, A4 => 
                           n15609, ZN => n15618);
   U13815 : AOI22_X1 port map( A1 => REGISTERS_28_44_port, A2 => n16570, B1 => 
                           REGISTERS_31_44_port, B2 => n16583, ZN => n15616);
   U13816 : AOI22_X1 port map( A1 => REGISTERS_26_44_port, A2 => n16582, B1 => 
                           REGISTERS_29_44_port, B2 => n16574, ZN => n15615);
   U13817 : AOI22_X1 port map( A1 => REGISTERS_10_44_port, A2 => n16560, B1 => 
                           REGISTERS_16_44_port, B2 => n16561, ZN => n15614);
   U13818 : AOI22_X1 port map( A1 => REGISTERS_9_44_port, A2 => n16029, B1 => 
                           REGISTERS_22_44_port, B2 => n16556, ZN => n15613);
   U13819 : NAND4_X1 port map( A1 => n15616, A2 => n15615, A3 => n15614, A4 => 
                           n15613, ZN => n15617);
   U13820 : NOR3_X1 port map( A1 => n15619, A2 => n15618, A3 => n15617, ZN => 
                           n15625);
   U13821 : AOI22_X1 port map( A1 => REGISTERS_4_44_port, A2 => n16595, B1 => 
                           REGISTERS_6_44_port, B2 => n16546, ZN => n15623);
   U13822 : AOI22_X1 port map( A1 => REGISTERS_5_44_port, A2 => n16518, B1 => 
                           REGISTERS_0_44_port, B2 => n16547, ZN => n15622);
   U13823 : AOI22_X1 port map( A1 => REGISTERS_2_44_port, A2 => n16545, B1 => 
                           REGISTERS_1_44_port, B2 => n16544, ZN => n15621);
   U13824 : AOI22_X1 port map( A1 => REGISTERS_7_44_port, A2 => n16454, B1 => 
                           REGISTERS_3_44_port, B2 => n16593, ZN => n15620);
   U13825 : AND4_X1 port map( A1 => n15623, A2 => n15622, A3 => n15621, A4 => 
                           n15620, ZN => n15624);
   U13826 : OAI222_X1 port map( A1 => n15796, A2 => n15625, B1 => n16553, B2 =>
                           n15624, C1 => n16026, C2 => n8422, ZN => n8589);
   U13827 : AOI22_X1 port map( A1 => REGISTERS_18_43_port, A2 => n16584, B1 => 
                           REGISTERS_12_43_port, B2 => n16580, ZN => n15629);
   U13828 : AOI22_X1 port map( A1 => REGISTERS_17_43_port, A2 => n16579, B1 => 
                           REGISTERS_29_43_port, B2 => n16574, ZN => n15628);
   U13829 : AOI22_X1 port map( A1 => REGISTERS_24_43_port, A2 => n16559, B1 => 
                           REGISTERS_21_43_port, B2 => n16568, ZN => n15627);
   U13830 : AOI22_X1 port map( A1 => REGISTERS_11_43_port, A2 => n16414, B1 => 
                           REGISTERS_28_43_port, B2 => n16570, ZN => n15626);
   U13831 : NAND4_X1 port map( A1 => n15629, A2 => n15628, A3 => n15627, A4 => 
                           n15626, ZN => n15640);
   U13832 : AOI22_X1 port map( A1 => REGISTERS_30_43_port, A2 => n16555, B1 => 
                           REGISTERS_14_43_port, B2 => n16571, ZN => n15633);
   U13833 : AOI22_X1 port map( A1 => REGISTERS_19_43_port, A2 => n16569, B1 => 
                           REGISTERS_22_43_port, B2 => n16556, ZN => n15632);
   U13834 : AOI22_X1 port map( A1 => REGISTERS_16_43_port, A2 => n16561, B1 => 
                           REGISTERS_27_43_port, B2 => n16573, ZN => n15631);
   U13835 : AOI22_X1 port map( A1 => REGISTERS_20_43_port, A2 => n16581, B1 => 
                           REGISTERS_13_43_port, B2 => n16562, ZN => n15630);
   U13836 : NAND4_X1 port map( A1 => n15633, A2 => n15632, A3 => n15631, A4 => 
                           n15630, ZN => n15639);
   U13837 : AOI22_X1 port map( A1 => REGISTERS_15_43_port, A2 => n16558, B1 => 
                           REGISTERS_8_43_port, B2 => n16567, ZN => n15637);
   U13838 : AOI22_X1 port map( A1 => REGISTERS_23_43_port, A2 => n16572, B1 => 
                           REGISTERS_31_43_port, B2 => n16583, ZN => n15636);
   U13839 : AOI22_X1 port map( A1 => REGISTERS_10_43_port, A2 => n16560, B1 => 
                           REGISTERS_26_43_port, B2 => n16582, ZN => n15635);
   U13840 : AOI22_X1 port map( A1 => REGISTERS_9_43_port, A2 => n16029, B1 => 
                           REGISTERS_25_43_port, B2 => n16557, ZN => n15634);
   U13841 : NAND4_X1 port map( A1 => n15637, A2 => n15636, A3 => n15635, A4 => 
                           n15634, ZN => n15638);
   U13842 : NOR3_X1 port map( A1 => n15640, A2 => n15639, A3 => n15638, ZN => 
                           n15646);
   U13843 : AOI22_X1 port map( A1 => REGISTERS_6_43_port, A2 => n16592, B1 => 
                           REGISTERS_1_43_port, B2 => n16544, ZN => n15644);
   U13844 : AOI22_X1 port map( A1 => REGISTERS_0_43_port, A2 => n16547, B1 => 
                           REGISTERS_3_43_port, B2 => n16453, ZN => n15643);
   U13845 : AOI22_X1 port map( A1 => REGISTERS_5_43_port, A2 => n16215, B1 => 
                           REGISTERS_4_43_port, B2 => n16595, ZN => n15642);
   U13846 : AOI22_X1 port map( A1 => REGISTERS_2_43_port, A2 => n16545, B1 => 
                           REGISTERS_7_43_port, B2 => n16594, ZN => n15641);
   U13847 : AND4_X1 port map( A1 => n15644, A2 => n15643, A3 => n15642, A4 => 
                           n15641, ZN => n15645);
   U13848 : OAI222_X1 port map( A1 => n15796, A2 => n15646, B1 => n16553, B2 =>
                           n15645, C1 => n16049, C2 => n8421, ZN => n8590);
   U13849 : AOI22_X1 port map( A1 => REGISTERS_16_42_port, A2 => n16561, B1 => 
                           REGISTERS_11_42_port, B2 => n15782, ZN => n15650);
   U13850 : AOI22_X1 port map( A1 => REGISTERS_8_42_port, A2 => n16567, B1 => 
                           REGISTERS_17_42_port, B2 => n16579, ZN => n15649);
   U13851 : AOI22_X1 port map( A1 => REGISTERS_19_42_port, A2 => n16569, B1 => 
                           REGISTERS_9_42_port, B2 => n16029, ZN => n15648);
   U13852 : AOI22_X1 port map( A1 => REGISTERS_27_42_port, A2 => n16573, B1 => 
                           REGISTERS_15_42_port, B2 => n16558, ZN => n15647);
   U13853 : NAND4_X1 port map( A1 => n15650, A2 => n15649, A3 => n15648, A4 => 
                           n15647, ZN => n15661);
   U13854 : AOI22_X1 port map( A1 => REGISTERS_13_42_port, A2 => n16562, B1 => 
                           REGISTERS_25_42_port, B2 => n16557, ZN => n15654);
   U13855 : AOI22_X1 port map( A1 => REGISTERS_26_42_port, A2 => n16582, B1 => 
                           REGISTERS_18_42_port, B2 => n16584, ZN => n15653);
   U13856 : AOI22_X1 port map( A1 => REGISTERS_30_42_port, A2 => n16555, B1 => 
                           REGISTERS_14_42_port, B2 => n16571, ZN => n15652);
   U13857 : AOI22_X1 port map( A1 => REGISTERS_21_42_port, A2 => n16568, B1 => 
                           REGISTERS_29_42_port, B2 => n16574, ZN => n15651);
   U13858 : NAND4_X1 port map( A1 => n15654, A2 => n15653, A3 => n15652, A4 => 
                           n15651, ZN => n15660);
   U13859 : AOI22_X1 port map( A1 => REGISTERS_10_42_port, A2 => n16560, B1 => 
                           REGISTERS_12_42_port, B2 => n16580, ZN => n15658);
   U13860 : AOI22_X1 port map( A1 => REGISTERS_22_42_port, A2 => n16556, B1 => 
                           REGISTERS_24_42_port, B2 => n16559, ZN => n15657);
   U13861 : AOI22_X1 port map( A1 => REGISTERS_23_42_port, A2 => n16572, B1 => 
                           REGISTERS_20_42_port, B2 => n16581, ZN => n15656);
   U13862 : AOI22_X1 port map( A1 => REGISTERS_31_42_port, A2 => n16583, B1 => 
                           REGISTERS_28_42_port, B2 => n16570, ZN => n15655);
   U13863 : NAND4_X1 port map( A1 => n15658, A2 => n15657, A3 => n15656, A4 => 
                           n15655, ZN => n15659);
   U13864 : NOR3_X1 port map( A1 => n15661, A2 => n15660, A3 => n15659, ZN => 
                           n15667);
   U13865 : AOI22_X1 port map( A1 => REGISTERS_7_42_port, A2 => n16594, B1 => 
                           REGISTERS_0_42_port, B2 => n16547, ZN => n15665);
   U13866 : AOI22_X1 port map( A1 => REGISTERS_1_42_port, A2 => n16544, B1 => 
                           REGISTERS_4_42_port, B2 => n16543, ZN => n15664);
   U13867 : AOI22_X1 port map( A1 => REGISTERS_3_42_port, A2 => n15746, B1 => 
                           REGISTERS_6_42_port, B2 => n16546, ZN => n15663);
   U13868 : AOI22_X1 port map( A1 => REGISTERS_5_42_port, A2 => n16215, B1 => 
                           REGISTERS_2_42_port, B2 => n16596, ZN => n15662);
   U13869 : OAI222_X1 port map( A1 => n15796, A2 => n15667, B1 => n16553, B2 =>
                           n15666, C1 => n16026, C2 => n8420, ZN => n8591);
   U13870 : AOI22_X1 port map( A1 => REGISTERS_22_41_port, A2 => n16556, B1 => 
                           REGISTERS_29_41_port, B2 => n16574, ZN => n15671);
   U13871 : AOI22_X1 port map( A1 => REGISTERS_18_41_port, A2 => n16584, B1 => 
                           REGISTERS_28_41_port, B2 => n16570, ZN => n15670);
   U13872 : AOI22_X1 port map( A1 => REGISTERS_9_41_port, A2 => n16029, B1 => 
                           REGISTERS_15_41_port, B2 => n16558, ZN => n15669);
   U13873 : AOI22_X1 port map( A1 => REGISTERS_30_41_port, A2 => n16555, B1 => 
                           REGISTERS_13_41_port, B2 => n16562, ZN => n15668);
   U13874 : NAND4_X1 port map( A1 => n15671, A2 => n15670, A3 => n15669, A4 => 
                           n15668, ZN => n15682);
   U13875 : AOI22_X1 port map( A1 => REGISTERS_12_41_port, A2 => n16580, B1 => 
                           REGISTERS_25_41_port, B2 => n16557, ZN => n15675);
   U13876 : AOI22_X1 port map( A1 => REGISTERS_10_41_port, A2 => n16560, B1 => 
                           REGISTERS_26_41_port, B2 => n16582, ZN => n15674);
   U13877 : AOI22_X1 port map( A1 => REGISTERS_23_41_port, A2 => n16572, B1 => 
                           REGISTERS_20_41_port, B2 => n16581, ZN => n15673);
   U13878 : AOI22_X1 port map( A1 => REGISTERS_14_41_port, A2 => n16571, B1 => 
                           REGISTERS_24_41_port, B2 => n16559, ZN => n15672);
   U13879 : NAND4_X1 port map( A1 => n15675, A2 => n15674, A3 => n15673, A4 => 
                           n15672, ZN => n15681);
   U13880 : AOI22_X1 port map( A1 => REGISTERS_27_41_port, A2 => n16573, B1 => 
                           REGISTERS_21_41_port, B2 => n16568, ZN => n15679);
   U13881 : AOI22_X1 port map( A1 => REGISTERS_8_41_port, A2 => n16567, B1 => 
                           REGISTERS_31_41_port, B2 => n16583, ZN => n15678);
   U13882 : AOI22_X1 port map( A1 => REGISTERS_16_41_port, A2 => n16561, B1 => 
                           REGISTERS_17_41_port, B2 => n16579, ZN => n15677);
   U13883 : AOI22_X1 port map( A1 => REGISTERS_11_41_port, A2 => n15782, B1 => 
                           REGISTERS_19_41_port, B2 => n16569, ZN => n15676);
   U13884 : NAND4_X1 port map( A1 => n15679, A2 => n15678, A3 => n15677, A4 => 
                           n15676, ZN => n15680);
   U13885 : NOR3_X1 port map( A1 => n15682, A2 => n15681, A3 => n15680, ZN => 
                           n15688);
   U13886 : AOI22_X1 port map( A1 => REGISTERS_4_41_port, A2 => n16543, B1 => 
                           REGISTERS_0_41_port, B2 => n16597, ZN => n15686);
   U13887 : AOI22_X1 port map( A1 => REGISTERS_5_41_port, A2 => n16215, B1 => 
                           REGISTERS_2_41_port, B2 => n16545, ZN => n15685);
   U13888 : AOI22_X1 port map( A1 => REGISTERS_3_41_port, A2 => n16453, B1 => 
                           REGISTERS_6_41_port, B2 => n16546, ZN => n15684);
   U13889 : AOI22_X1 port map( A1 => REGISTERS_7_41_port, A2 => n16216, B1 => 
                           REGISTERS_1_41_port, B2 => n16544, ZN => n15683);
   U13890 : AND4_X1 port map( A1 => n15686, A2 => n15685, A3 => n15684, A4 => 
                           n15683, ZN => n15687);
   U13891 : OAI222_X1 port map( A1 => n15796, A2 => n15688, B1 => n16553, B2 =>
                           n15687, C1 => n16049, C2 => n8419, ZN => n8592);
   U13892 : AOI22_X1 port map( A1 => REGISTERS_14_40_port, A2 => n16571, B1 => 
                           REGISTERS_19_40_port, B2 => n16569, ZN => n15692);
   U13893 : AOI22_X1 port map( A1 => REGISTERS_24_40_port, A2 => n16559, B1 => 
                           REGISTERS_12_40_port, B2 => n16580, ZN => n15691);
   U13894 : AOI22_X1 port map( A1 => REGISTERS_29_40_port, A2 => n16574, B1 => 
                           REGISTERS_23_40_port, B2 => n16572, ZN => n15690);
   U13895 : AOI22_X1 port map( A1 => REGISTERS_15_40_port, A2 => n16558, B1 => 
                           REGISTERS_26_40_port, B2 => n16582, ZN => n15689);
   U13896 : NAND4_X1 port map( A1 => n15692, A2 => n15691, A3 => n15690, A4 => 
                           n15689, ZN => n15703);
   U13897 : AOI22_X1 port map( A1 => REGISTERS_9_40_port, A2 => n16029, B1 => 
                           REGISTERS_25_40_port, B2 => n16557, ZN => n15696);
   U13898 : AOI22_X1 port map( A1 => REGISTERS_13_40_port, A2 => n16562, B1 => 
                           REGISTERS_10_40_port, B2 => n16560, ZN => n15695);
   U13899 : AOI22_X1 port map( A1 => REGISTERS_21_40_port, A2 => n16568, B1 => 
                           REGISTERS_18_40_port, B2 => n16584, ZN => n15694);
   U13900 : AOI22_X1 port map( A1 => REGISTERS_20_40_port, A2 => n16581, B1 => 
                           REGISTERS_17_40_port, B2 => n16579, ZN => n15693);
   U13901 : NAND4_X1 port map( A1 => n15696, A2 => n15695, A3 => n15694, A4 => 
                           n15693, ZN => n15702);
   U13902 : AOI22_X1 port map( A1 => REGISTERS_27_40_port, A2 => n16573, B1 => 
                           REGISTERS_8_40_port, B2 => n16567, ZN => n15700);
   U13903 : AOI22_X1 port map( A1 => REGISTERS_31_40_port, A2 => n16583, B1 => 
                           REGISTERS_16_40_port, B2 => n16561, ZN => n15699);
   U13904 : AOI22_X1 port map( A1 => REGISTERS_30_40_port, A2 => n16555, B1 => 
                           REGISTERS_11_40_port, B2 => n15782, ZN => n15698);
   U13905 : AOI22_X1 port map( A1 => REGISTERS_22_40_port, A2 => n16556, B1 => 
                           REGISTERS_28_40_port, B2 => n16570, ZN => n15697);
   U13906 : NAND4_X1 port map( A1 => n15700, A2 => n15699, A3 => n15698, A4 => 
                           n15697, ZN => n15701);
   U13907 : NOR3_X1 port map( A1 => n15703, A2 => n15702, A3 => n15701, ZN => 
                           n15709);
   U13908 : AOI22_X1 port map( A1 => REGISTERS_6_40_port, A2 => n16546, B1 => 
                           REGISTERS_3_40_port, B2 => n16453, ZN => n15707);
   U13909 : AOI22_X1 port map( A1 => REGISTERS_5_40_port, A2 => n16215, B1 => 
                           REGISTERS_0_40_port, B2 => n16547, ZN => n15706);
   U13910 : AOI22_X1 port map( A1 => REGISTERS_7_40_port, A2 => n16216, B1 => 
                           REGISTERS_4_40_port, B2 => n16595, ZN => n15705);
   U13911 : AOI22_X1 port map( A1 => REGISTERS_2_40_port, A2 => n16545, B1 => 
                           REGISTERS_1_40_port, B2 => n16544, ZN => n15704);
   U13912 : AND4_X1 port map( A1 => n15707, A2 => n15706, A3 => n15705, A4 => 
                           n15704, ZN => n15708);
   U13913 : OAI222_X1 port map( A1 => n15796, A2 => n15709, B1 => n16553, B2 =>
                           n15708, C1 => n16026, C2 => n8418, ZN => n8593);
   U13914 : AOI22_X1 port map( A1 => REGISTERS_24_39_port, A2 => n16559, B1 => 
                           REGISTERS_13_39_port, B2 => n16562, ZN => n15713);
   U13915 : AOI22_X1 port map( A1 => REGISTERS_8_39_port, A2 => n16567, B1 => 
                           REGISTERS_17_39_port, B2 => n16579, ZN => n15712);
   U13916 : AOI22_X1 port map( A1 => REGISTERS_19_39_port, A2 => n16569, B1 => 
                           REGISTERS_28_39_port, B2 => n16570, ZN => n15711);
   U13917 : AOI22_X1 port map( A1 => REGISTERS_18_39_port, A2 => n16584, B1 => 
                           REGISTERS_29_39_port, B2 => n16574, ZN => n15710);
   U13918 : NAND4_X1 port map( A1 => n15713, A2 => n15712, A3 => n15711, A4 => 
                           n15710, ZN => n15724);
   U13919 : AOI22_X1 port map( A1 => REGISTERS_31_39_port, A2 => n16583, B1 => 
                           REGISTERS_20_39_port, B2 => n16581, ZN => n15717);
   U13920 : AOI22_X1 port map( A1 => REGISTERS_21_39_port, A2 => n16568, B1 => 
                           REGISTERS_26_39_port, B2 => n16582, ZN => n15716);
   U13921 : AOI22_X1 port map( A1 => REGISTERS_23_39_port, A2 => n16572, B1 => 
                           REGISTERS_25_39_port, B2 => n16557, ZN => n15715);
   U13922 : AOI22_X1 port map( A1 => REGISTERS_27_39_port, A2 => n16573, B1 => 
                           REGISTERS_14_39_port, B2 => n16571, ZN => n15714);
   U13923 : NAND4_X1 port map( A1 => n15717, A2 => n15716, A3 => n15715, A4 => 
                           n15714, ZN => n15723);
   U13924 : AOI22_X1 port map( A1 => REGISTERS_15_39_port, A2 => n16558, B1 => 
                           REGISTERS_16_39_port, B2 => n16561, ZN => n15721);
   U13925 : AOI22_X1 port map( A1 => REGISTERS_9_39_port, A2 => n16437, B1 => 
                           REGISTERS_10_39_port, B2 => n16560, ZN => n15720);
   U13926 : AOI22_X1 port map( A1 => REGISTERS_30_39_port, A2 => n16555, B1 => 
                           REGISTERS_22_39_port, B2 => n16556, ZN => n15719);
   U13927 : AOI22_X1 port map( A1 => REGISTERS_11_39_port, A2 => n16414, B1 => 
                           REGISTERS_12_39_port, B2 => n16580, ZN => n15718);
   U13928 : NAND4_X1 port map( A1 => n15721, A2 => n15720, A3 => n15719, A4 => 
                           n15718, ZN => n15722);
   U13929 : NOR3_X1 port map( A1 => n15724, A2 => n15723, A3 => n15722, ZN => 
                           n15730);
   U13930 : AOI22_X1 port map( A1 => REGISTERS_4_39_port, A2 => n16543, B1 => 
                           REGISTERS_3_39_port, B2 => n16593, ZN => n15728);
   U13931 : AOI22_X1 port map( A1 => REGISTERS_2_39_port, A2 => n16545, B1 => 
                           REGISTERS_1_39_port, B2 => n16544, ZN => n15727);
   U13932 : AOI22_X1 port map( A1 => REGISTERS_7_39_port, A2 => n16216, B1 => 
                           REGISTERS_0_39_port, B2 => n16547, ZN => n15726);
   U13933 : AOI22_X1 port map( A1 => REGISTERS_5_39_port, A2 => n16542, B1 => 
                           REGISTERS_6_39_port, B2 => n16546, ZN => n15725);
   U13934 : AND4_X1 port map( A1 => n15728, A2 => n15727, A3 => n15726, A4 => 
                           n15725, ZN => n15729);
   U13935 : OAI222_X1 port map( A1 => n15796, A2 => n15730, B1 => n16553, B2 =>
                           n15729, C1 => n16049, C2 => n8417, ZN => n8594);
   U13936 : AOI22_X1 port map( A1 => REGISTERS_16_38_port, A2 => n16561, B1 => 
                           REGISTERS_12_38_port, B2 => n16580, ZN => n15734);
   U13937 : AOI22_X1 port map( A1 => REGISTERS_18_38_port, A2 => n16584, B1 => 
                           REGISTERS_15_38_port, B2 => n16558, ZN => n15733);
   U13938 : AOI22_X1 port map( A1 => REGISTERS_30_38_port, A2 => n16555, B1 => 
                           REGISTERS_31_38_port, B2 => n16583, ZN => n15732);
   U13939 : AOI22_X1 port map( A1 => REGISTERS_11_38_port, A2 => n15782, B1 => 
                           REGISTERS_9_38_port, B2 => n16029, ZN => n15731);
   U13940 : NAND4_X1 port map( A1 => n15734, A2 => n15733, A3 => n15732, A4 => 
                           n15731, ZN => n15745);
   U13941 : AOI22_X1 port map( A1 => REGISTERS_25_38_port, A2 => n16557, B1 => 
                           REGISTERS_20_38_port, B2 => n16581, ZN => n15738);
   U13942 : AOI22_X1 port map( A1 => REGISTERS_29_38_port, A2 => n16574, B1 => 
                           REGISTERS_23_38_port, B2 => n16572, ZN => n15737);
   U13943 : AOI22_X1 port map( A1 => REGISTERS_8_38_port, A2 => n16567, B1 => 
                           REGISTERS_21_38_port, B2 => n16568, ZN => n15736);
   U13944 : AOI22_X1 port map( A1 => REGISTERS_28_38_port, A2 => n16570, B1 => 
                           REGISTERS_14_38_port, B2 => n16571, ZN => n15735);
   U13945 : NAND4_X1 port map( A1 => n15738, A2 => n15737, A3 => n15736, A4 => 
                           n15735, ZN => n15744);
   U13946 : AOI22_X1 port map( A1 => REGISTERS_13_38_port, A2 => n16562, B1 => 
                           REGISTERS_27_38_port, B2 => n16573, ZN => n15742);
   U13947 : AOI22_X1 port map( A1 => REGISTERS_24_38_port, A2 => n16559, B1 => 
                           REGISTERS_19_38_port, B2 => n16569, ZN => n15741);
   U13948 : AOI22_X1 port map( A1 => REGISTERS_26_38_port, A2 => n16582, B1 => 
                           REGISTERS_22_38_port, B2 => n16556, ZN => n15740);
   U13949 : AOI22_X1 port map( A1 => REGISTERS_10_38_port, A2 => n16560, B1 => 
                           REGISTERS_17_38_port, B2 => n16579, ZN => n15739);
   U13950 : NAND4_X1 port map( A1 => n15742, A2 => n15741, A3 => n15740, A4 => 
                           n15739, ZN => n15743);
   U13951 : NOR3_X1 port map( A1 => n15745, A2 => n15744, A3 => n15743, ZN => 
                           n15752);
   U13952 : AOI22_X1 port map( A1 => REGISTERS_5_38_port, A2 => n16518, B1 => 
                           REGISTERS_6_38_port, B2 => n16546, ZN => n15750);
   U13953 : AOI22_X1 port map( A1 => REGISTERS_2_38_port, A2 => n16545, B1 => 
                           REGISTERS_7_38_port, B2 => n16454, ZN => n15749);
   U13954 : AOI22_X1 port map( A1 => REGISTERS_3_38_port, A2 => n15746, B1 => 
                           REGISTERS_0_38_port, B2 => n16547, ZN => n15748);
   U13955 : AOI22_X1 port map( A1 => REGISTERS_4_38_port, A2 => n16595, B1 => 
                           REGISTERS_1_38_port, B2 => n16430, ZN => n15747);
   U13956 : AND4_X1 port map( A1 => n15750, A2 => n15749, A3 => n15748, A4 => 
                           n15747, ZN => n15751);
   U13957 : OAI222_X1 port map( A1 => n15796, A2 => n15752, B1 => n16553, B2 =>
                           n15751, C1 => n16026, C2 => n8416, ZN => n8595);
   U13958 : AOI22_X1 port map( A1 => REGISTERS_23_37_port, A2 => n16572, B1 => 
                           REGISTERS_29_37_port, B2 => n16574, ZN => n15756);
   U13959 : AOI22_X1 port map( A1 => REGISTERS_15_37_port, A2 => n16558, B1 => 
                           REGISTERS_11_37_port, B2 => n15782, ZN => n15755);
   U13960 : AOI22_X1 port map( A1 => REGISTERS_17_37_port, A2 => n16579, B1 => 
                           REGISTERS_30_37_port, B2 => n16555, ZN => n15754);
   U13961 : AOI22_X1 port map( A1 => REGISTERS_16_37_port, A2 => n16561, B1 => 
                           REGISTERS_21_37_port, B2 => n16568, ZN => n15753);
   U13962 : NAND4_X1 port map( A1 => n15756, A2 => n15755, A3 => n15754, A4 => 
                           n15753, ZN => n15767);
   U13963 : AOI22_X1 port map( A1 => REGISTERS_27_37_port, A2 => n16573, B1 => 
                           REGISTERS_8_37_port, B2 => n16567, ZN => n15760);
   U13964 : AOI22_X1 port map( A1 => REGISTERS_26_37_port, A2 => n16582, B1 => 
                           REGISTERS_22_37_port, B2 => n16556, ZN => n15759);
   U13965 : AOI22_X1 port map( A1 => REGISTERS_20_37_port, A2 => n16581, B1 => 
                           REGISTERS_18_37_port, B2 => n16584, ZN => n15758);
   U13966 : AOI22_X1 port map( A1 => REGISTERS_10_37_port, A2 => n16560, B1 => 
                           REGISTERS_24_37_port, B2 => n16559, ZN => n15757);
   U13967 : NAND4_X1 port map( A1 => n15760, A2 => n15759, A3 => n15758, A4 => 
                           n15757, ZN => n15766);
   U13968 : AOI22_X1 port map( A1 => REGISTERS_28_37_port, A2 => n16570, B1 => 
                           REGISTERS_31_37_port, B2 => n16583, ZN => n15764);
   U13969 : AOI22_X1 port map( A1 => REGISTERS_19_37_port, A2 => n16569, B1 => 
                           REGISTERS_25_37_port, B2 => n16557, ZN => n15763);
   U13970 : AOI22_X1 port map( A1 => REGISTERS_12_37_port, A2 => n16580, B1 => 
                           REGISTERS_13_37_port, B2 => n16562, ZN => n15762);
   U13971 : AOI22_X1 port map( A1 => REGISTERS_9_37_port, A2 => n16437, B1 => 
                           REGISTERS_14_37_port, B2 => n16571, ZN => n15761);
   U13972 : NAND4_X1 port map( A1 => n15764, A2 => n15763, A3 => n15762, A4 => 
                           n15761, ZN => n15765);
   U13973 : NOR3_X1 port map( A1 => n15767, A2 => n15766, A3 => n15765, ZN => 
                           n15773);
   U13974 : AOI22_X1 port map( A1 => REGISTERS_4_37_port, A2 => n16543, B1 => 
                           REGISTERS_5_37_port, B2 => n16518, ZN => n15771);
   U13975 : AOI22_X1 port map( A1 => REGISTERS_6_37_port, A2 => n16592, B1 => 
                           REGISTERS_7_37_port, B2 => n16594, ZN => n15770);
   U13976 : AOI22_X1 port map( A1 => REGISTERS_2_37_port, A2 => n16545, B1 => 
                           REGISTERS_0_37_port, B2 => n16597, ZN => n15769);
   U13977 : AOI22_X1 port map( A1 => REGISTERS_3_37_port, A2 => n16453, B1 => 
                           REGISTERS_1_37_port, B2 => n16544, ZN => n15768);
   U13978 : AND4_X1 port map( A1 => n15771, A2 => n15770, A3 => n15769, A4 => 
                           n15768, ZN => n15772);
   U13979 : OAI222_X1 port map( A1 => n15796, A2 => n15773, B1 => n16553, B2 =>
                           n15772, C1 => n16049, C2 => n8415, ZN => n8596);
   U13980 : AOI22_X1 port map( A1 => REGISTERS_28_36_port, A2 => n16570, B1 => 
                           REGISTERS_16_36_port, B2 => n16561, ZN => n15777);
   U13981 : AOI22_X1 port map( A1 => REGISTERS_26_36_port, A2 => n16582, B1 => 
                           REGISTERS_9_36_port, B2 => n16029, ZN => n15776);
   U13982 : AOI22_X1 port map( A1 => REGISTERS_18_36_port, A2 => n16584, B1 => 
                           REGISTERS_27_36_port, B2 => n16573, ZN => n15775);
   U13983 : AOI22_X1 port map( A1 => REGISTERS_31_36_port, A2 => n16583, B1 => 
                           REGISTERS_17_36_port, B2 => n16579, ZN => n15774);
   U13984 : NAND4_X1 port map( A1 => n15777, A2 => n15776, A3 => n15775, A4 => 
                           n15774, ZN => n15789);
   U13985 : AOI22_X1 port map( A1 => REGISTERS_30_36_port, A2 => n16555, B1 => 
                           REGISTERS_13_36_port, B2 => n16562, ZN => n15781);
   U13986 : AOI22_X1 port map( A1 => REGISTERS_29_36_port, A2 => n16574, B1 => 
                           REGISTERS_12_36_port, B2 => n16580, ZN => n15780);
   U13987 : AOI22_X1 port map( A1 => REGISTERS_22_36_port, A2 => n16556, B1 => 
                           REGISTERS_24_36_port, B2 => n16559, ZN => n15779);
   U13988 : AOI22_X1 port map( A1 => REGISTERS_23_36_port, A2 => n16572, B1 => 
                           REGISTERS_15_36_port, B2 => n16558, ZN => n15778);
   U13989 : NAND4_X1 port map( A1 => n15781, A2 => n15780, A3 => n15779, A4 => 
                           n15778, ZN => n15788);
   U13990 : AOI22_X1 port map( A1 => REGISTERS_8_36_port, A2 => n16567, B1 => 
                           REGISTERS_14_36_port, B2 => n16571, ZN => n15786);
   U13991 : AOI22_X1 port map( A1 => REGISTERS_19_36_port, A2 => n16569, B1 => 
                           REGISTERS_20_36_port, B2 => n16581, ZN => n15785);
   U13992 : AOI22_X1 port map( A1 => REGISTERS_25_36_port, A2 => n16557, B1 => 
                           REGISTERS_21_36_port, B2 => n16568, ZN => n15784);
   U13993 : AOI22_X1 port map( A1 => REGISTERS_10_36_port, A2 => n16560, B1 => 
                           REGISTERS_11_36_port, B2 => n15782, ZN => n15783);
   U13994 : NAND4_X1 port map( A1 => n15786, A2 => n15785, A3 => n15784, A4 => 
                           n15783, ZN => n15787);
   U13995 : NOR3_X1 port map( A1 => n15789, A2 => n15788, A3 => n15787, ZN => 
                           n15795);
   U13996 : AOI22_X1 port map( A1 => REGISTERS_3_36_port, A2 => n16453, B1 => 
                           REGISTERS_6_36_port, B2 => n16546, ZN => n15793);
   U13997 : AOI22_X1 port map( A1 => REGISTERS_0_36_port, A2 => n16547, B1 => 
                           REGISTERS_1_36_port, B2 => n16430, ZN => n15792);
   U13998 : AOI22_X1 port map( A1 => REGISTERS_7_36_port, A2 => n16216, B1 => 
                           REGISTERS_2_36_port, B2 => n16596, ZN => n15791);
   U13999 : AOI22_X1 port map( A1 => REGISTERS_5_36_port, A2 => n16542, B1 => 
                           REGISTERS_4_36_port, B2 => n16543, ZN => n15790);
   U14000 : AND4_X1 port map( A1 => n15793, A2 => n15792, A3 => n15791, A4 => 
                           n15790, ZN => n15794);
   U14001 : OAI222_X1 port map( A1 => n15796, A2 => n15795, B1 => n16553, B2 =>
                           n15794, C1 => n16026, C2 => n8414, ZN => n8597);
   U14002 : AOI22_X1 port map( A1 => REGISTERS_27_35_port, A2 => n16573, B1 => 
                           REGISTERS_8_35_port, B2 => n16567, ZN => n15800);
   U14003 : AOI22_X1 port map( A1 => REGISTERS_13_35_port, A2 => n16562, B1 => 
                           REGISTERS_11_35_port, B2 => n15782, ZN => n15799);
   U14004 : AOI22_X1 port map( A1 => REGISTERS_12_35_port, A2 => n16580, B1 => 
                           REGISTERS_17_35_port, B2 => n16579, ZN => n15798);
   U14005 : AOI22_X1 port map( A1 => REGISTERS_22_35_port, A2 => n16556, B1 => 
                           REGISTERS_28_35_port, B2 => n16570, ZN => n15797);
   U14006 : NAND4_X1 port map( A1 => n15800, A2 => n15799, A3 => n15798, A4 => 
                           n15797, ZN => n15811);
   U14007 : AOI22_X1 port map( A1 => REGISTERS_26_35_port, A2 => n16582, B1 => 
                           REGISTERS_19_35_port, B2 => n16569, ZN => n15804);
   U14008 : AOI22_X1 port map( A1 => REGISTERS_21_35_port, A2 => n16568, B1 => 
                           REGISTERS_15_35_port, B2 => n16558, ZN => n15803);
   U14009 : AOI22_X1 port map( A1 => REGISTERS_29_35_port, A2 => n16574, B1 => 
                           REGISTERS_16_35_port, B2 => n16561, ZN => n15802);
   U14010 : AOI22_X1 port map( A1 => REGISTERS_20_35_port, A2 => n16581, B1 => 
                           REGISTERS_24_35_port, B2 => n16559, ZN => n15801);
   U14011 : NAND4_X1 port map( A1 => n15804, A2 => n15803, A3 => n15802, A4 => 
                           n15801, ZN => n15810);
   U14012 : AOI22_X1 port map( A1 => REGISTERS_18_35_port, A2 => n16584, B1 => 
                           REGISTERS_9_35_port, B2 => n16029, ZN => n15808);
   U14013 : AOI22_X1 port map( A1 => REGISTERS_23_35_port, A2 => n16572, B1 => 
                           REGISTERS_14_35_port, B2 => n16571, ZN => n15807);
   U14014 : AOI22_X1 port map( A1 => REGISTERS_30_35_port, A2 => n16555, B1 => 
                           REGISTERS_31_35_port, B2 => n16583, ZN => n15806);
   U14015 : AOI22_X1 port map( A1 => REGISTERS_25_35_port, A2 => n16557, B1 => 
                           REGISTERS_10_35_port, B2 => n16560, ZN => n15805);
   U14016 : NAND4_X1 port map( A1 => n15808, A2 => n15807, A3 => n15806, A4 => 
                           n15805, ZN => n15809);
   U14017 : NOR3_X1 port map( A1 => n15811, A2 => n15810, A3 => n15809, ZN => 
                           n15817);
   U14018 : AOI22_X1 port map( A1 => REGISTERS_1_35_port, A2 => n16322, B1 => 
                           REGISTERS_6_35_port, B2 => n16546, ZN => n15815);
   U14019 : AOI22_X1 port map( A1 => REGISTERS_5_35_port, A2 => n16542, B1 => 
                           REGISTERS_0_35_port, B2 => n16547, ZN => n15814);
   U14020 : AOI22_X1 port map( A1 => REGISTERS_4_35_port, A2 => n16543, B1 => 
                           REGISTERS_7_35_port, B2 => n16594, ZN => n15813);
   U14021 : AOI22_X1 port map( A1 => REGISTERS_3_35_port, A2 => n16593, B1 => 
                           REGISTERS_2_35_port, B2 => n16545, ZN => n15812);
   U14022 : OAI222_X1 port map( A1 => n15796, A2 => n15817, B1 => n16553, B2 =>
                           n15816, C1 => n16026, C2 => n8413, ZN => n8598);
   U14023 : AOI22_X1 port map( A1 => REGISTERS_26_34_port, A2 => n16582, B1 => 
                           REGISTERS_25_34_port, B2 => n16557, ZN => n15821);
   U14024 : AOI22_X1 port map( A1 => REGISTERS_28_34_port, A2 => n16570, B1 => 
                           REGISTERS_8_34_port, B2 => n16567, ZN => n15820);
   U14025 : AOI22_X1 port map( A1 => REGISTERS_9_34_port, A2 => n16525, B1 => 
                           REGISTERS_31_34_port, B2 => n16583, ZN => n15819);
   U14026 : AOI22_X1 port map( A1 => REGISTERS_21_34_port, A2 => n16568, B1 => 
                           REGISTERS_17_34_port, B2 => n16579, ZN => n15818);
   U14027 : NAND4_X1 port map( A1 => n15821, A2 => n15820, A3 => n15819, A4 => 
                           n15818, ZN => n15832);
   U14028 : AOI22_X1 port map( A1 => REGISTERS_11_34_port, A2 => n16530, B1 => 
                           REGISTERS_20_34_port, B2 => n16581, ZN => n15825);
   U14029 : AOI22_X1 port map( A1 => REGISTERS_30_34_port, A2 => n16555, B1 => 
                           REGISTERS_27_34_port, B2 => n16573, ZN => n15824);
   U14030 : AOI22_X1 port map( A1 => REGISTERS_12_34_port, A2 => n16580, B1 => 
                           REGISTERS_16_34_port, B2 => n16561, ZN => n15823);
   U14031 : AOI22_X1 port map( A1 => REGISTERS_14_34_port, A2 => n16571, B1 => 
                           REGISTERS_18_34_port, B2 => n16584, ZN => n15822);
   U14032 : NAND4_X1 port map( A1 => n15825, A2 => n15824, A3 => n15823, A4 => 
                           n15822, ZN => n15831);
   U14033 : AOI22_X1 port map( A1 => REGISTERS_13_34_port, A2 => n16562, B1 => 
                           REGISTERS_22_34_port, B2 => n16556, ZN => n15829);
   U14034 : AOI22_X1 port map( A1 => REGISTERS_24_34_port, A2 => n16559, B1 => 
                           REGISTERS_23_34_port, B2 => n16572, ZN => n15828);
   U14035 : AOI22_X1 port map( A1 => REGISTERS_19_34_port, A2 => n16569, B1 => 
                           REGISTERS_15_34_port, B2 => n16558, ZN => n15827);
   U14036 : AOI22_X1 port map( A1 => REGISTERS_29_34_port, A2 => n16574, B1 => 
                           REGISTERS_10_34_port, B2 => n16560, ZN => n15826);
   U14037 : NAND4_X1 port map( A1 => n15829, A2 => n15828, A3 => n15827, A4 => 
                           n15826, ZN => n15830);
   U14038 : NOR3_X1 port map( A1 => n15832, A2 => n15831, A3 => n15830, ZN => 
                           n15838);
   U14039 : AOI22_X1 port map( A1 => REGISTERS_7_34_port, A2 => n16454, B1 => 
                           REGISTERS_1_34_port, B2 => n16430, ZN => n15836);
   U14040 : AOI22_X1 port map( A1 => REGISTERS_6_34_port, A2 => n16592, B1 => 
                           REGISTERS_3_34_port, B2 => n16593, ZN => n15835);
   U14041 : AOI22_X1 port map( A1 => REGISTERS_0_34_port, A2 => n16547, B1 => 
                           REGISTERS_5_34_port, B2 => n16542, ZN => n15834);
   U14042 : AOI22_X1 port map( A1 => REGISTERS_2_34_port, A2 => n16545, B1 => 
                           REGISTERS_4_34_port, B2 => n16543, ZN => n15833);
   U14043 : AND4_X1 port map( A1 => n15836, A2 => n15835, A3 => n15834, A4 => 
                           n15833, ZN => n15837);
   U14044 : OAI222_X1 port map( A1 => n15796, A2 => n15838, B1 => n16553, B2 =>
                           n15837, C1 => n16049, C2 => n8412, ZN => n8599);
   U14045 : AOI22_X1 port map( A1 => REGISTERS_23_33_port, A2 => n16572, B1 => 
                           REGISTERS_26_33_port, B2 => n16582, ZN => n15842);
   U14046 : AOI22_X1 port map( A1 => REGISTERS_11_33_port, A2 => n16530, B1 => 
                           REGISTERS_13_33_port, B2 => n16562, ZN => n15841);
   U14047 : AOI22_X1 port map( A1 => REGISTERS_24_33_port, A2 => n16559, B1 => 
                           REGISTERS_18_33_port, B2 => n16584, ZN => n15840);
   U14048 : AOI22_X1 port map( A1 => REGISTERS_28_33_port, A2 => n16570, B1 => 
                           REGISTERS_19_33_port, B2 => n16569, ZN => n15839);
   U14049 : NAND4_X1 port map( A1 => n15842, A2 => n15841, A3 => n15840, A4 => 
                           n15839, ZN => n15853);
   U14050 : AOI22_X1 port map( A1 => REGISTERS_21_33_port, A2 => n16568, B1 => 
                           REGISTERS_22_33_port, B2 => n16556, ZN => n15846);
   U14051 : AOI22_X1 port map( A1 => REGISTERS_14_33_port, A2 => n16571, B1 => 
                           REGISTERS_25_33_port, B2 => n16557, ZN => n15845);
   U14052 : AOI22_X1 port map( A1 => REGISTERS_9_33_port, A2 => n16525, B1 => 
                           REGISTERS_8_33_port, B2 => n16567, ZN => n15844);
   U14053 : AOI22_X1 port map( A1 => REGISTERS_10_33_port, A2 => n16560, B1 => 
                           REGISTERS_16_33_port, B2 => n16561, ZN => n15843);
   U14054 : NAND4_X1 port map( A1 => n15846, A2 => n15845, A3 => n15844, A4 => 
                           n15843, ZN => n15852);
   U14055 : AOI22_X1 port map( A1 => REGISTERS_12_33_port, A2 => n16580, B1 => 
                           REGISTERS_27_33_port, B2 => n16573, ZN => n15850);
   U14056 : AOI22_X1 port map( A1 => REGISTERS_20_33_port, A2 => n16581, B1 => 
                           REGISTERS_31_33_port, B2 => n16583, ZN => n15849);
   U14057 : AOI22_X1 port map( A1 => REGISTERS_29_33_port, A2 => n16574, B1 => 
                           REGISTERS_17_33_port, B2 => n16579, ZN => n15848);
   U14058 : AOI22_X1 port map( A1 => REGISTERS_15_33_port, A2 => n16558, B1 => 
                           REGISTERS_30_33_port, B2 => n16555, ZN => n15847);
   U14059 : NAND4_X1 port map( A1 => n15850, A2 => n15849, A3 => n15848, A4 => 
                           n15847, ZN => n15851);
   U14060 : NOR3_X1 port map( A1 => n15853, A2 => n15852, A3 => n15851, ZN => 
                           n15859);
   U14061 : AOI22_X1 port map( A1 => REGISTERS_2_33_port, A2 => n16545, B1 => 
                           REGISTERS_3_33_port, B2 => n16593, ZN => n15857);
   U14062 : AOI22_X1 port map( A1 => REGISTERS_7_33_port, A2 => n16594, B1 => 
                           REGISTERS_1_33_port, B2 => n16430, ZN => n15856);
   U14063 : AOI22_X1 port map( A1 => REGISTERS_5_33_port, A2 => n16518, B1 => 
                           REGISTERS_0_33_port, B2 => n16547, ZN => n15855);
   U14064 : AOI22_X1 port map( A1 => REGISTERS_6_33_port, A2 => n16592, B1 => 
                           REGISTERS_4_33_port, B2 => n16595, ZN => n15854);
   U14065 : AND4_X1 port map( A1 => n15857, A2 => n15856, A3 => n15855, A4 => 
                           n15854, ZN => n15858);
   U14066 : OAI222_X1 port map( A1 => n16605, A2 => n15859, B1 => n16553, B2 =>
                           n15858, C1 => n16026, C2 => n8411, ZN => n8600);
   U14067 : AOI22_X1 port map( A1 => REGISTERS_24_32_port, A2 => n16559, B1 => 
                           REGISTERS_20_32_port, B2 => n16581, ZN => n15863);
   U14068 : AOI22_X1 port map( A1 => REGISTERS_22_32_port, A2 => n16556, B1 => 
                           REGISTERS_19_32_port, B2 => n16569, ZN => n15862);
   U14069 : AOI22_X1 port map( A1 => REGISTERS_18_32_port, A2 => n16584, B1 => 
                           REGISTERS_31_32_port, B2 => n16583, ZN => n15861);
   U14070 : AOI22_X1 port map( A1 => REGISTERS_16_32_port, A2 => n16561, B1 => 
                           REGISTERS_14_32_port, B2 => n16571, ZN => n15860);
   U14071 : NAND4_X1 port map( A1 => n15863, A2 => n15862, A3 => n15861, A4 => 
                           n15860, ZN => n15874);
   U14072 : AOI22_X1 port map( A1 => REGISTERS_17_32_port, A2 => n16579, B1 => 
                           REGISTERS_30_32_port, B2 => n16555, ZN => n15867);
   U14073 : AOI22_X1 port map( A1 => REGISTERS_27_32_port, A2 => n16573, B1 => 
                           REGISTERS_25_32_port, B2 => n16557, ZN => n15866);
   U14074 : AOI22_X1 port map( A1 => REGISTERS_9_32_port, A2 => n16029, B1 => 
                           REGISTERS_26_32_port, B2 => n16582, ZN => n15865);
   U14075 : AOI22_X1 port map( A1 => REGISTERS_15_32_port, A2 => n16558, B1 => 
                           REGISTERS_12_32_port, B2 => n16580, ZN => n15864);
   U14076 : NAND4_X1 port map( A1 => n15867, A2 => n15866, A3 => n15865, A4 => 
                           n15864, ZN => n15873);
   U14077 : AOI22_X1 port map( A1 => REGISTERS_28_32_port, A2 => n16570, B1 => 
                           REGISTERS_29_32_port, B2 => n16574, ZN => n15871);
   U14078 : AOI22_X1 port map( A1 => REGISTERS_21_32_port, A2 => n16568, B1 => 
                           REGISTERS_11_32_port, B2 => n16414, ZN => n15870);
   U14079 : AOI22_X1 port map( A1 => REGISTERS_10_32_port, A2 => n16560, B1 => 
                           REGISTERS_8_32_port, B2 => n16567, ZN => n15869);
   U14080 : AOI22_X1 port map( A1 => REGISTERS_13_32_port, A2 => n16562, B1 => 
                           REGISTERS_23_32_port, B2 => n16572, ZN => n15868);
   U14081 : NAND4_X1 port map( A1 => n15871, A2 => n15870, A3 => n15869, A4 => 
                           n15868, ZN => n15872);
   U14082 : NOR3_X1 port map( A1 => n15874, A2 => n15873, A3 => n15872, ZN => 
                           n15880);
   U14083 : AOI22_X1 port map( A1 => REGISTERS_3_32_port, A2 => n16593, B1 => 
                           REGISTERS_1_32_port, B2 => n16430, ZN => n15878);
   U14084 : AOI22_X1 port map( A1 => REGISTERS_4_32_port, A2 => n16595, B1 => 
                           REGISTERS_0_32_port, B2 => n16547, ZN => n15877);
   U14085 : AOI22_X1 port map( A1 => REGISTERS_7_32_port, A2 => n16454, B1 => 
                           REGISTERS_6_32_port, B2 => n16546, ZN => n15876);
   U14086 : AOI22_X1 port map( A1 => REGISTERS_5_32_port, A2 => n16518, B1 => 
                           REGISTERS_2_32_port, B2 => n16596, ZN => n15875);
   U14087 : AND4_X1 port map( A1 => n15878, A2 => n15877, A3 => n15876, A4 => 
                           n15875, ZN => n15879);
   U14088 : OAI222_X1 port map( A1 => n15796, A2 => n15880, B1 => n16553, B2 =>
                           n15879, C1 => n16049, C2 => n8410, ZN => n8601);
   U14089 : AOI22_X1 port map( A1 => REGISTERS_11_31_port, A2 => n16530, B1 => 
                           REGISTERS_8_31_port, B2 => n16567, ZN => n15884);
   U14090 : AOI22_X1 port map( A1 => REGISTERS_15_31_port, A2 => n16558, B1 => 
                           REGISTERS_21_31_port, B2 => n16568, ZN => n15883);
   U14091 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n16581, B1 => 
                           REGISTERS_18_31_port, B2 => n16584, ZN => n15882);
   U14092 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n16556, B1 => 
                           REGISTERS_13_31_port, B2 => n16562, ZN => n15881);
   U14093 : NAND4_X1 port map( A1 => n15884, A2 => n15883, A3 => n15882, A4 => 
                           n15881, ZN => n15895);
   U14094 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n16525, B1 => 
                           REGISTERS_12_31_port, B2 => n16580, ZN => n15888);
   U14095 : AOI22_X1 port map( A1 => REGISTERS_27_31_port, A2 => n16573, B1 => 
                           REGISTERS_26_31_port, B2 => n16582, ZN => n15887);
   U14096 : AOI22_X1 port map( A1 => REGISTERS_19_31_port, A2 => n16569, B1 => 
                           REGISTERS_30_31_port, B2 => n16555, ZN => n15886);
   U14097 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n16574, B1 => 
                           REGISTERS_24_31_port, B2 => n16559, ZN => n15885);
   U14098 : NAND4_X1 port map( A1 => n15888, A2 => n15887, A3 => n15886, A4 => 
                           n15885, ZN => n15894);
   U14099 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n16570, B1 => 
                           REGISTERS_10_31_port, B2 => n16560, ZN => n15892);
   U14100 : AOI22_X1 port map( A1 => REGISTERS_23_31_port, A2 => n16572, B1 => 
                           REGISTERS_31_31_port, B2 => n16583, ZN => n15891);
   U14101 : AOI22_X1 port map( A1 => REGISTERS_14_31_port, A2 => n16571, B1 => 
                           REGISTERS_25_31_port, B2 => n16557, ZN => n15890);
   U14102 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n16561, B1 => 
                           REGISTERS_17_31_port, B2 => n16579, ZN => n15889);
   U14103 : NAND4_X1 port map( A1 => n15892, A2 => n15891, A3 => n15890, A4 => 
                           n15889, ZN => n15893);
   U14104 : NOR3_X1 port map( A1 => n15895, A2 => n15894, A3 => n15893, ZN => 
                           n15901);
   U14105 : AOI22_X1 port map( A1 => REGISTERS_0_31_port, A2 => n16597, B1 => 
                           REGISTERS_2_31_port, B2 => n16545, ZN => n15899);
   U14106 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n16543, B1 => 
                           REGISTERS_3_31_port, B2 => n16593, ZN => n15898);
   U14107 : AOI22_X1 port map( A1 => REGISTERS_7_31_port, A2 => n16594, B1 => 
                           REGISTERS_6_31_port, B2 => n16546, ZN => n15897);
   U14108 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n16542, B1 => 
                           REGISTERS_1_31_port, B2 => n16430, ZN => n15896);
   U14109 : AND4_X1 port map( A1 => n15899, A2 => n15898, A3 => n15897, A4 => 
                           n15896, ZN => n15900);
   U14110 : OAI222_X1 port map( A1 => n15796, A2 => n15901, B1 => n16553, B2 =>
                           n15900, C1 => n16026, C2 => n8409, ZN => n8602);
   U14111 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n16570, B1 => 
                           REGISTERS_9_30_port, B2 => n16029, ZN => n15905);
   U14112 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n16579, B1 => 
                           REGISTERS_27_30_port, B2 => n16573, ZN => n15904);
   U14113 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n16581, B1 => 
                           REGISTERS_14_30_port, B2 => n16571, ZN => n15903);
   U14114 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n16557, B1 => 
                           REGISTERS_16_30_port, B2 => n16561, ZN => n15902);
   U14115 : NAND4_X1 port map( A1 => n15905, A2 => n15904, A3 => n15903, A4 => 
                           n15902, ZN => n15916);
   U14116 : AOI22_X1 port map( A1 => REGISTERS_15_30_port, A2 => n16558, B1 => 
                           REGISTERS_24_30_port, B2 => n16559, ZN => n15909);
   U14117 : AOI22_X1 port map( A1 => REGISTERS_18_30_port, A2 => n16584, B1 => 
                           REGISTERS_31_30_port, B2 => n16583, ZN => n15908);
   U14118 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n16562, B1 => 
                           REGISTERS_12_30_port, B2 => n16580, ZN => n15907);
   U14119 : AOI22_X1 port map( A1 => REGISTERS_22_30_port, A2 => n16556, B1 => 
                           REGISTERS_21_30_port, B2 => n16568, ZN => n15906);
   U14120 : NAND4_X1 port map( A1 => n15909, A2 => n15908, A3 => n15907, A4 => 
                           n15906, ZN => n15915);
   U14121 : AOI22_X1 port map( A1 => REGISTERS_23_30_port, A2 => n16572, B1 => 
                           REGISTERS_11_30_port, B2 => n15782, ZN => n15913);
   U14122 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n16567, B1 => 
                           REGISTERS_19_30_port, B2 => n16569, ZN => n15912);
   U14123 : AOI22_X1 port map( A1 => REGISTERS_10_30_port, A2 => n16560, B1 => 
                           REGISTERS_26_30_port, B2 => n16582, ZN => n15911);
   U14124 : AOI22_X1 port map( A1 => REGISTERS_30_30_port, A2 => n16555, B1 => 
                           REGISTERS_29_30_port, B2 => n16574, ZN => n15910);
   U14125 : NAND4_X1 port map( A1 => n15913, A2 => n15912, A3 => n15911, A4 => 
                           n15910, ZN => n15914);
   U14126 : NOR3_X1 port map( A1 => n15916, A2 => n15915, A3 => n15914, ZN => 
                           n15922);
   U14127 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n16544, B1 => 
                           REGISTERS_7_30_port, B2 => n16594, ZN => n15920);
   U14128 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n16542, B1 => 
                           REGISTERS_2_30_port, B2 => n16596, ZN => n15919);
   U14129 : AOI22_X1 port map( A1 => REGISTERS_0_30_port, A2 => n16597, B1 => 
                           REGISTERS_4_30_port, B2 => n16543, ZN => n15918);
   U14130 : AOI22_X1 port map( A1 => REGISTERS_3_30_port, A2 => n16453, B1 => 
                           REGISTERS_6_30_port, B2 => n16546, ZN => n15917);
   U14131 : AND4_X1 port map( A1 => n15920, A2 => n15919, A3 => n15918, A4 => 
                           n15917, ZN => n15921);
   U14132 : OAI222_X1 port map( A1 => n16605, A2 => n15922, B1 => n16553, B2 =>
                           n15921, C1 => n16049, C2 => n8408, ZN => n8603);
   U14133 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n16579, B1 => 
                           REGISTERS_19_29_port, B2 => n16569, ZN => n15926);
   U14134 : AOI22_X1 port map( A1 => REGISTERS_31_29_port, A2 => n16583, B1 => 
                           REGISTERS_8_29_port, B2 => n16567, ZN => n15925);
   U14135 : AOI22_X1 port map( A1 => REGISTERS_14_29_port, A2 => n16571, B1 => 
                           REGISTERS_28_29_port, B2 => n16570, ZN => n15924);
   U14136 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n16559, B1 => 
                           REGISTERS_27_29_port, B2 => n16573, ZN => n15923);
   U14137 : NAND4_X1 port map( A1 => n15926, A2 => n15925, A3 => n15924, A4 => 
                           n15923, ZN => n15937);
   U14138 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n16557, B1 => 
                           REGISTERS_22_29_port, B2 => n16556, ZN => n15930);
   U14139 : AOI22_X1 port map( A1 => REGISTERS_26_29_port, A2 => n16582, B1 => 
                           REGISTERS_20_29_port, B2 => n16581, ZN => n15929);
   U14140 : AOI22_X1 port map( A1 => REGISTERS_15_29_port, A2 => n16558, B1 => 
                           REGISTERS_9_29_port, B2 => n16029, ZN => n15928);
   U14141 : AOI22_X1 port map( A1 => REGISTERS_30_29_port, A2 => n16555, B1 => 
                           REGISTERS_13_29_port, B2 => n16562, ZN => n15927);
   U14142 : NAND4_X1 port map( A1 => n15930, A2 => n15929, A3 => n15928, A4 => 
                           n15927, ZN => n15936);
   U14143 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n16580, B1 => 
                           REGISTERS_23_29_port, B2 => n16572, ZN => n15934);
   U14144 : AOI22_X1 port map( A1 => REGISTERS_11_29_port, A2 => n15782, B1 => 
                           REGISTERS_21_29_port, B2 => n16568, ZN => n15933);
   U14145 : AOI22_X1 port map( A1 => REGISTERS_18_29_port, A2 => n16584, B1 => 
                           REGISTERS_16_29_port, B2 => n16561, ZN => n15932);
   U14146 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n16574, B1 => 
                           REGISTERS_10_29_port, B2 => n16560, ZN => n15931);
   U14147 : NAND4_X1 port map( A1 => n15934, A2 => n15933, A3 => n15932, A4 => 
                           n15931, ZN => n15935);
   U14148 : NOR3_X1 port map( A1 => n15937, A2 => n15936, A3 => n15935, ZN => 
                           n15943);
   U14149 : AOI22_X1 port map( A1 => REGISTERS_7_29_port, A2 => n16594, B1 => 
                           REGISTERS_4_29_port, B2 => n16595, ZN => n15941);
   U14150 : AOI22_X1 port map( A1 => REGISTERS_3_29_port, A2 => n16593, B1 => 
                           REGISTERS_1_29_port, B2 => n16430, ZN => n15940);
   U14151 : AOI22_X1 port map( A1 => REGISTERS_6_29_port, A2 => n16592, B1 => 
                           REGISTERS_2_29_port, B2 => n16596, ZN => n15939);
   U14152 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n16547, B1 => 
                           REGISTERS_5_29_port, B2 => n16518, ZN => n15938);
   U14153 : AND4_X1 port map( A1 => n15941, A2 => n15940, A3 => n15939, A4 => 
                           n15938, ZN => n15942);
   U14154 : OAI222_X1 port map( A1 => n16605, A2 => n15943, B1 => n16553, B2 =>
                           n15942, C1 => n16026, C2 => n8407, ZN => n8604);
   U14155 : AOI22_X1 port map( A1 => REGISTERS_30_28_port, A2 => n16555, B1 => 
                           REGISTERS_12_28_port, B2 => n16580, ZN => n15947);
   U14156 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n16437, B1 => 
                           REGISTERS_21_28_port, B2 => n16568, ZN => n15946);
   U14157 : AOI22_X1 port map( A1 => REGISTERS_10_28_port, A2 => n16560, B1 => 
                           REGISTERS_13_28_port, B2 => n16562, ZN => n15945);
   U14158 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n16557, B1 => 
                           REGISTERS_29_28_port, B2 => n16574, ZN => n15944);
   U14159 : NAND4_X1 port map( A1 => n15947, A2 => n15946, A3 => n15945, A4 => 
                           n15944, ZN => n15958);
   U14160 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n16579, B1 => 
                           REGISTERS_27_28_port, B2 => n16573, ZN => n15951);
   U14161 : AOI22_X1 port map( A1 => REGISTERS_15_28_port, A2 => n16558, B1 => 
                           REGISTERS_24_28_port, B2 => n16559, ZN => n15950);
   U14162 : AOI22_X1 port map( A1 => REGISTERS_14_28_port, A2 => n16571, B1 => 
                           REGISTERS_8_28_port, B2 => n16567, ZN => n15949);
   U14163 : AOI22_X1 port map( A1 => REGISTERS_26_28_port, A2 => n16582, B1 => 
                           REGISTERS_19_28_port, B2 => n16569, ZN => n15948);
   U14164 : NAND4_X1 port map( A1 => n15951, A2 => n15950, A3 => n15949, A4 => 
                           n15948, ZN => n15957);
   U14165 : AOI22_X1 port map( A1 => REGISTERS_18_28_port, A2 => n16584, B1 => 
                           REGISTERS_28_28_port, B2 => n16570, ZN => n15955);
   U14166 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n16581, B1 => 
                           REGISTERS_23_28_port, B2 => n16572, ZN => n15954);
   U14167 : AOI22_X1 port map( A1 => REGISTERS_22_28_port, A2 => n16556, B1 => 
                           REGISTERS_11_28_port, B2 => n16414, ZN => n15953);
   U14168 : AOI22_X1 port map( A1 => REGISTERS_31_28_port, A2 => n16583, B1 => 
                           REGISTERS_16_28_port, B2 => n16561, ZN => n15952);
   U14169 : NAND4_X1 port map( A1 => n15955, A2 => n15954, A3 => n15953, A4 => 
                           n15952, ZN => n15956);
   U14170 : NOR3_X1 port map( A1 => n15958, A2 => n15957, A3 => n15956, ZN => 
                           n15964);
   U14171 : AOI22_X1 port map( A1 => REGISTERS_6_28_port, A2 => n16344, B1 => 
                           REGISTERS_2_28_port, B2 => n16545, ZN => n15962);
   U14172 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n16543, B1 => 
                           REGISTERS_1_28_port, B2 => n16430, ZN => n15961);
   U14173 : AOI22_X1 port map( A1 => REGISTERS_3_28_port, A2 => n16453, B1 => 
                           REGISTERS_7_28_port, B2 => n16594, ZN => n15960);
   U14174 : AOI22_X1 port map( A1 => REGISTERS_0_28_port, A2 => n16547, B1 => 
                           REGISTERS_5_28_port, B2 => n16518, ZN => n15959);
   U14175 : AND4_X1 port map( A1 => n15962, A2 => n15961, A3 => n15960, A4 => 
                           n15959, ZN => n15963);
   U14176 : OAI222_X1 port map( A1 => n15796, A2 => n15964, B1 => n16553, B2 =>
                           n15963, C1 => n16049, C2 => n8406, ZN => n8605);
   U14177 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n16574, B1 => 
                           REGISTERS_17_27_port, B2 => n16579, ZN => n15968);
   U14178 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n16567, B1 => 
                           REGISTERS_23_27_port, B2 => n16572, ZN => n15967);
   U14179 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n16580, B1 => 
                           REGISTERS_30_27_port, B2 => n16555, ZN => n15966);
   U14180 : AOI22_X1 port map( A1 => REGISTERS_27_27_port, A2 => n16573, B1 => 
                           REGISTERS_10_27_port, B2 => n16560, ZN => n15965);
   U14181 : NAND4_X1 port map( A1 => n15968, A2 => n15967, A3 => n15966, A4 => 
                           n15965, ZN => n15979);
   U14182 : AOI22_X1 port map( A1 => REGISTERS_15_27_port, A2 => n16558, B1 => 
                           REGISTERS_20_27_port, B2 => n16581, ZN => n15972);
   U14183 : AOI22_X1 port map( A1 => REGISTERS_14_27_port, A2 => n16571, B1 => 
                           REGISTERS_18_27_port, B2 => n16584, ZN => n15971);
   U14184 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n16568, B1 => 
                           REGISTERS_22_27_port, B2 => n16556, ZN => n15970);
   U14185 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n16525, B1 => 
                           REGISTERS_11_27_port, B2 => n15782, ZN => n15969);
   U14186 : NAND4_X1 port map( A1 => n15972, A2 => n15971, A3 => n15970, A4 => 
                           n15969, ZN => n15978);
   U14187 : AOI22_X1 port map( A1 => REGISTERS_19_27_port, A2 => n16569, B1 => 
                           REGISTERS_16_27_port, B2 => n16561, ZN => n15976);
   U14188 : AOI22_X1 port map( A1 => REGISTERS_31_27_port, A2 => n16583, B1 => 
                           REGISTERS_13_27_port, B2 => n16562, ZN => n15975);
   U14189 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n16557, B1 => 
                           REGISTERS_26_27_port, B2 => n16582, ZN => n15974);
   U14190 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n16570, B1 => 
                           REGISTERS_24_27_port, B2 => n16559, ZN => n15973);
   U14191 : NAND4_X1 port map( A1 => n15976, A2 => n15975, A3 => n15974, A4 => 
                           n15973, ZN => n15977);
   U14192 : NOR3_X1 port map( A1 => n15979, A2 => n15978, A3 => n15977, ZN => 
                           n15985);
   U14193 : AOI22_X1 port map( A1 => REGISTERS_2_27_port, A2 => n16545, B1 => 
                           REGISTERS_4_27_port, B2 => n16543, ZN => n15983);
   U14194 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n16430, B1 => 
                           REGISTERS_5_27_port, B2 => n16518, ZN => n15982);
   U14195 : AOI22_X1 port map( A1 => REGISTERS_6_27_port, A2 => n16592, B1 => 
                           REGISTERS_3_27_port, B2 => n16593, ZN => n15981);
   U14196 : AOI22_X1 port map( A1 => REGISTERS_7_27_port, A2 => n16454, B1 => 
                           REGISTERS_0_27_port, B2 => n16547, ZN => n15980);
   U14197 : AND4_X1 port map( A1 => n15983, A2 => n15982, A3 => n15981, A4 => 
                           n15980, ZN => n15984);
   U14198 : OAI222_X1 port map( A1 => n16605, A2 => n15985, B1 => n16603, B2 =>
                           n15984, C1 => n16026, C2 => n8405, ZN => n8606);
   U14199 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n16557, B1 => 
                           REGISTERS_15_26_port, B2 => n16558, ZN => n15989);
   U14200 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n16562, B1 => 
                           REGISTERS_17_26_port, B2 => n16579, ZN => n15988);
   U14201 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n16525, B1 => 
                           REGISTERS_14_26_port, B2 => n16571, ZN => n15987);
   U14202 : AOI22_X1 port map( A1 => REGISTERS_27_26_port, A2 => n16573, B1 => 
                           REGISTERS_21_26_port, B2 => n16568, ZN => n15986);
   U14203 : NAND4_X1 port map( A1 => n15989, A2 => n15988, A3 => n15987, A4 => 
                           n15986, ZN => n16000);
   U14204 : AOI22_X1 port map( A1 => REGISTERS_23_26_port, A2 => n16572, B1 => 
                           REGISTERS_28_26_port, B2 => n16570, ZN => n15993);
   U14205 : AOI22_X1 port map( A1 => REGISTERS_31_26_port, A2 => n16583, B1 => 
                           REGISTERS_22_26_port, B2 => n16556, ZN => n15992);
   U14206 : AOI22_X1 port map( A1 => REGISTERS_11_26_port, A2 => n16414, B1 => 
                           REGISTERS_12_26_port, B2 => n16580, ZN => n15991);
   U14207 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n16574, B1 => 
                           REGISTERS_20_26_port, B2 => n16581, ZN => n15990);
   U14208 : NAND4_X1 port map( A1 => n15993, A2 => n15992, A3 => n15991, A4 => 
                           n15990, ZN => n15999);
   U14209 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n16567, B1 => 
                           REGISTERS_10_26_port, B2 => n16560, ZN => n15997);
   U14210 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n16559, B1 => 
                           REGISTERS_18_26_port, B2 => n16584, ZN => n15996);
   U14211 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n16561, B1 => 
                           REGISTERS_30_26_port, B2 => n16555, ZN => n15995);
   U14212 : AOI22_X1 port map( A1 => REGISTERS_26_26_port, A2 => n16582, B1 => 
                           REGISTERS_19_26_port, B2 => n16569, ZN => n15994);
   U14213 : NAND4_X1 port map( A1 => n15997, A2 => n15996, A3 => n15995, A4 => 
                           n15994, ZN => n15998);
   U14214 : NOR3_X1 port map( A1 => n16000, A2 => n15999, A3 => n15998, ZN => 
                           n16006);
   U14215 : AOI22_X1 port map( A1 => REGISTERS_0_26_port, A2 => n16597, B1 => 
                           REGISTERS_5_26_port, B2 => n16518, ZN => n16004);
   U14216 : AOI22_X1 port map( A1 => REGISTERS_3_26_port, A2 => n16453, B1 => 
                           REGISTERS_7_26_port, B2 => n16594, ZN => n16003);
   U14217 : AOI22_X1 port map( A1 => REGISTERS_2_26_port, A2 => n16545, B1 => 
                           REGISTERS_6_26_port, B2 => n16546, ZN => n16002);
   U14218 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n16595, B1 => 
                           REGISTERS_1_26_port, B2 => n16430, ZN => n16001);
   U14219 : AND4_X1 port map( A1 => n16004, A2 => n16003, A3 => n16002, A4 => 
                           n16001, ZN => n16005);
   U14220 : OAI222_X1 port map( A1 => n15796, A2 => n16006, B1 => n16603, B2 =>
                           n16005, C1 => n16049, C2 => n8404, ZN => n8607);
   U14221 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n16568, B1 => 
                           REGISTERS_16_25_port, B2 => n16561, ZN => n16010);
   U14222 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n16581, B1 => 
                           REGISTERS_11_25_port, B2 => n16414, ZN => n16009);
   U14223 : AOI22_X1 port map( A1 => REGISTERS_14_25_port, A2 => n16571, B1 => 
                           REGISTERS_28_25_port, B2 => n16570, ZN => n16008);
   U14224 : AOI22_X1 port map( A1 => REGISTERS_26_25_port, A2 => n16582, B1 => 
                           REGISTERS_25_25_port, B2 => n16557, ZN => n16007);
   U14225 : NAND4_X1 port map( A1 => n16010, A2 => n16009, A3 => n16008, A4 => 
                           n16007, ZN => n16021);
   U14226 : AOI22_X1 port map( A1 => REGISTERS_30_25_port, A2 => n16555, B1 => 
                           REGISTERS_15_25_port, B2 => n16558, ZN => n16014);
   U14227 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n16567, B1 => 
                           REGISTERS_9_25_port, B2 => n16029, ZN => n16013);
   U14228 : AOI22_X1 port map( A1 => REGISTERS_18_25_port, A2 => n16584, B1 => 
                           REGISTERS_13_25_port, B2 => n16562, ZN => n16012);
   U14229 : AOI22_X1 port map( A1 => REGISTERS_10_25_port, A2 => n16560, B1 => 
                           REGISTERS_23_25_port, B2 => n16572, ZN => n16011);
   U14230 : NAND4_X1 port map( A1 => n16014, A2 => n16013, A3 => n16012, A4 => 
                           n16011, ZN => n16020);
   U14231 : AOI22_X1 port map( A1 => REGISTERS_22_25_port, A2 => n16556, B1 => 
                           REGISTERS_29_25_port, B2 => n16574, ZN => n16018);
   U14232 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n16559, B1 => 
                           REGISTERS_31_25_port, B2 => n16583, ZN => n16017);
   U14233 : AOI22_X1 port map( A1 => REGISTERS_27_25_port, A2 => n16573, B1 => 
                           REGISTERS_12_25_port, B2 => n16580, ZN => n16016);
   U14234 : AOI22_X1 port map( A1 => REGISTERS_19_25_port, A2 => n16569, B1 => 
                           REGISTERS_17_25_port, B2 => n16579, ZN => n16015);
   U14235 : NAND4_X1 port map( A1 => n16018, A2 => n16017, A3 => n16016, A4 => 
                           n16015, ZN => n16019);
   U14236 : NOR3_X1 port map( A1 => n16021, A2 => n16020, A3 => n16019, ZN => 
                           n16028);
   U14237 : AOI22_X1 port map( A1 => REGISTERS_0_25_port, A2 => n16597, B1 => 
                           REGISTERS_4_25_port, B2 => n16595, ZN => n16025);
   U14238 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n16542, B1 => 
                           REGISTERS_2_25_port, B2 => n16545, ZN => n16024);
   U14239 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n16322, B1 => 
                           REGISTERS_3_25_port, B2 => n16593, ZN => n16023);
   U14240 : AOI22_X1 port map( A1 => REGISTERS_6_25_port, A2 => n16344, B1 => 
                           REGISTERS_7_25_port, B2 => n16594, ZN => n16022);
   U14241 : AND4_X1 port map( A1 => n16025, A2 => n16024, A3 => n16023, A4 => 
                           n16022, ZN => n16027);
   U14242 : OAI222_X1 port map( A1 => n16605, A2 => n16028, B1 => n16603, B2 =>
                           n16027, C1 => n16026, C2 => n8403, ZN => n8608);
   U14243 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n16570, B1 => 
                           REGISTERS_9_24_port, B2 => n16029, ZN => n16033);
   U14244 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n16561, B1 => 
                           REGISTERS_21_24_port, B2 => n16568, ZN => n16032);
   U14245 : AOI22_X1 port map( A1 => REGISTERS_11_24_port, A2 => n15782, B1 => 
                           REGISTERS_23_24_port, B2 => n16572, ZN => n16031);
   U14246 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n16574, B1 => 
                           REGISTERS_26_24_port, B2 => n16582, ZN => n16030);
   U14247 : NAND4_X1 port map( A1 => n16033, A2 => n16032, A3 => n16031, A4 => 
                           n16030, ZN => n16044);
   U14248 : AOI22_X1 port map( A1 => REGISTERS_18_24_port, A2 => n16584, B1 => 
                           REGISTERS_25_24_port, B2 => n16557, ZN => n16037);
   U14249 : AOI22_X1 port map( A1 => REGISTERS_22_24_port, A2 => n16556, B1 => 
                           REGISTERS_15_24_port, B2 => n16558, ZN => n16036);
   U14250 : AOI22_X1 port map( A1 => REGISTERS_30_24_port, A2 => n16555, B1 => 
                           REGISTERS_10_24_port, B2 => n16560, ZN => n16035);
   U14251 : AOI22_X1 port map( A1 => REGISTERS_27_24_port, A2 => n16573, B1 => 
                           REGISTERS_13_24_port, B2 => n16562, ZN => n16034);
   U14252 : NAND4_X1 port map( A1 => n16037, A2 => n16036, A3 => n16035, A4 => 
                           n16034, ZN => n16043);
   U14253 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n16581, B1 => 
                           REGISTERS_19_24_port, B2 => n16569, ZN => n16041);
   U14254 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n16559, B1 => 
                           REGISTERS_12_24_port, B2 => n16580, ZN => n16040);
   U14255 : AOI22_X1 port map( A1 => REGISTERS_31_24_port, A2 => n16583, B1 => 
                           REGISTERS_8_24_port, B2 => n16567, ZN => n16039);
   U14256 : AOI22_X1 port map( A1 => REGISTERS_14_24_port, A2 => n16571, B1 => 
                           REGISTERS_17_24_port, B2 => n16579, ZN => n16038);
   U14257 : NAND4_X1 port map( A1 => n16041, A2 => n16040, A3 => n16039, A4 => 
                           n16038, ZN => n16042);
   U14258 : NOR3_X1 port map( A1 => n16044, A2 => n16043, A3 => n16042, ZN => 
                           n16051);
   U14259 : AOI22_X1 port map( A1 => REGISTERS_6_24_port, A2 => n16592, B1 => 
                           REGISTERS_1_24_port, B2 => n16430, ZN => n16048);
   U14260 : AOI22_X1 port map( A1 => REGISTERS_0_24_port, A2 => n16547, B1 => 
                           REGISTERS_5_24_port, B2 => n16518, ZN => n16047);
   U14261 : AOI22_X1 port map( A1 => REGISTERS_3_24_port, A2 => n16593, B1 => 
                           REGISTERS_2_24_port, B2 => n16596, ZN => n16046);
   U14262 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n16595, B1 => 
                           REGISTERS_7_24_port, B2 => n16594, ZN => n16045);
   U14263 : AND4_X1 port map( A1 => n16048, A2 => n16047, A3 => n16046, A4 => 
                           n16045, ZN => n16050);
   U14264 : OAI222_X1 port map( A1 => n15796, A2 => n16051, B1 => n16603, B2 =>
                           n16050, C1 => n16049, C2 => n8402, ZN => n8609);
   U14265 : AOI22_X1 port map( A1 => REGISTERS_15_23_port, A2 => n16558, B1 => 
                           REGISTERS_26_23_port, B2 => n16582, ZN => n16055);
   U14266 : AOI22_X1 port map( A1 => REGISTERS_14_23_port, A2 => n16571, B1 => 
                           REGISTERS_18_23_port, B2 => n16584, ZN => n16054);
   U14267 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n16567, B1 => 
                           REGISTERS_9_23_port, B2 => n16525, ZN => n16053);
   U14268 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n16559, B1 => 
                           REGISTERS_21_23_port, B2 => n16568, ZN => n16052);
   U14269 : NAND4_X1 port map( A1 => n16055, A2 => n16054, A3 => n16053, A4 => 
                           n16052, ZN => n16066);
   U14270 : AOI22_X1 port map( A1 => REGISTERS_31_23_port, A2 => n16583, B1 => 
                           REGISTERS_13_23_port, B2 => n16562, ZN => n16059);
   U14271 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n16557, B1 => 
                           REGISTERS_22_23_port, B2 => n16556, ZN => n16058);
   U14272 : AOI22_X1 port map( A1 => REGISTERS_10_23_port, A2 => n16560, B1 => 
                           REGISTERS_20_23_port, B2 => n16581, ZN => n16057);
   U14273 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n16561, B1 => 
                           REGISTERS_19_23_port, B2 => n16569, ZN => n16056);
   U14274 : NAND4_X1 port map( A1 => n16059, A2 => n16058, A3 => n16057, A4 => 
                           n16056, ZN => n16065);
   U14275 : AOI22_X1 port map( A1 => REGISTERS_30_23_port, A2 => n16555, B1 => 
                           REGISTERS_27_23_port, B2 => n16573, ZN => n16063);
   U14276 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n16579, B1 => 
                           REGISTERS_29_23_port, B2 => n16574, ZN => n16062);
   U14277 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n16580, B1 => 
                           REGISTERS_23_23_port, B2 => n16572, ZN => n16061);
   U14278 : AOI22_X1 port map( A1 => REGISTERS_11_23_port, A2 => n16414, B1 => 
                           REGISTERS_28_23_port, B2 => n16570, ZN => n16060);
   U14279 : NAND4_X1 port map( A1 => n16063, A2 => n16062, A3 => n16061, A4 => 
                           n16060, ZN => n16064);
   U14280 : NOR3_X1 port map( A1 => n16066, A2 => n16065, A3 => n16064, ZN => 
                           n16073);
   U14281 : AOI22_X1 port map( A1 => REGISTERS_3_23_port, A2 => n16453, B1 => 
                           REGISTERS_5_23_port, B2 => n16518, ZN => n16070);
   U14282 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n16543, B1 => 
                           REGISTERS_2_23_port, B2 => n16596, ZN => n16069);
   U14283 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n16544, B1 => 
                           REGISTERS_7_23_port, B2 => n16594, ZN => n16068);
   U14284 : AOI22_X1 port map( A1 => REGISTERS_6_23_port, A2 => n16592, B1 => 
                           REGISTERS_0_23_port, B2 => n16547, ZN => n16067);
   U14285 : AND4_X1 port map( A1 => n16070, A2 => n16069, A3 => n16068, A4 => 
                           n16067, ZN => n16072);
   U14286 : OAI222_X1 port map( A1 => n15796, A2 => n16073, B1 => n16603, B2 =>
                           n16072, C1 => n16071, C2 => n8401, ZN => n8610);
   U14287 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n16580, B1 => 
                           REGISTERS_25_22_port, B2 => n16557, ZN => n16077);
   U14288 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n16574, B1 => 
                           REGISTERS_17_22_port, B2 => n16579, ZN => n16076);
   U14289 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n16562, B1 => 
                           REGISTERS_19_22_port, B2 => n16569, ZN => n16075);
   U14290 : AOI22_X1 port map( A1 => REGISTERS_10_22_port, A2 => n16560, B1 => 
                           REGISTERS_9_22_port, B2 => n16525, ZN => n16074);
   U14291 : NAND4_X1 port map( A1 => n16077, A2 => n16076, A3 => n16075, A4 => 
                           n16074, ZN => n16088);
   U14292 : AOI22_X1 port map( A1 => REGISTERS_23_22_port, A2 => n16572, B1 => 
                           REGISTERS_18_22_port, B2 => n16584, ZN => n16081);
   U14293 : AOI22_X1 port map( A1 => REGISTERS_26_22_port, A2 => n16582, B1 => 
                           REGISTERS_24_22_port, B2 => n16559, ZN => n16080);
   U14294 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n16567, B1 => 
                           REGISTERS_11_22_port, B2 => n16414, ZN => n16079);
   U14295 : AOI22_X1 port map( A1 => REGISTERS_15_22_port, A2 => n16558, B1 => 
                           REGISTERS_20_22_port, B2 => n16581, ZN => n16078);
   U14296 : NAND4_X1 port map( A1 => n16081, A2 => n16080, A3 => n16079, A4 => 
                           n16078, ZN => n16087);
   U14297 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n16570, B1 => 
                           REGISTERS_27_22_port, B2 => n16573, ZN => n16085);
   U14298 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n16561, B1 => 
                           REGISTERS_22_22_port, B2 => n16556, ZN => n16084);
   U14299 : AOI22_X1 port map( A1 => REGISTERS_14_22_port, A2 => n16571, B1 => 
                           REGISTERS_30_22_port, B2 => n16555, ZN => n16083);
   U14300 : AOI22_X1 port map( A1 => REGISTERS_31_22_port, A2 => n16583, B1 => 
                           REGISTERS_21_22_port, B2 => n16568, ZN => n16082);
   U14301 : NAND4_X1 port map( A1 => n16085, A2 => n16084, A3 => n16083, A4 => 
                           n16082, ZN => n16086);
   U14302 : NOR3_X1 port map( A1 => n16088, A2 => n16087, A3 => n16086, ZN => 
                           n16094);
   U14303 : AOI22_X1 port map( A1 => REGISTERS_7_22_port, A2 => n16454, B1 => 
                           REGISTERS_1_22_port, B2 => n16430, ZN => n16092);
   U14304 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n16542, B1 => 
                           REGISTERS_0_22_port, B2 => n16547, ZN => n16091);
   U14305 : AOI22_X1 port map( A1 => REGISTERS_2_22_port, A2 => n16545, B1 => 
                           REGISTERS_4_22_port, B2 => n16543, ZN => n16090);
   U14306 : AOI22_X1 port map( A1 => REGISTERS_3_22_port, A2 => n16593, B1 => 
                           REGISTERS_6_22_port, B2 => n16546, ZN => n16089);
   U14307 : AND4_X1 port map( A1 => n16092, A2 => n16091, A3 => n16090, A4 => 
                           n16089, ZN => n16093);
   U14308 : OAI222_X1 port map( A1 => n15796, A2 => n16094, B1 => n16603, B2 =>
                           n16093, C1 => n16071, C2 => n8400, ZN => n8611);
   U14309 : AOI22_X1 port map( A1 => REGISTERS_11_21_port, A2 => n15782, B1 => 
                           REGISTERS_27_21_port, B2 => n16573, ZN => n16098);
   U14310 : AOI22_X1 port map( A1 => REGISTERS_18_21_port, A2 => n16584, B1 => 
                           REGISTERS_17_21_port, B2 => n16579, ZN => n16097);
   U14311 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n16581, B1 => 
                           REGISTERS_31_21_port, B2 => n16583, ZN => n16096);
   U14312 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n16568, B1 => 
                           REGISTERS_30_21_port, B2 => n16555, ZN => n16095);
   U14313 : NAND4_X1 port map( A1 => n16098, A2 => n16097, A3 => n16096, A4 => 
                           n16095, ZN => n16109);
   U14314 : AOI22_X1 port map( A1 => REGISTERS_10_21_port, A2 => n16560, B1 => 
                           REGISTERS_13_21_port, B2 => n16562, ZN => n16102);
   U14315 : AOI22_X1 port map( A1 => REGISTERS_26_21_port, A2 => n16582, B1 => 
                           REGISTERS_16_21_port, B2 => n16561, ZN => n16101);
   U14316 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n16525, B1 => 
                           REGISTERS_14_21_port, B2 => n16571, ZN => n16100);
   U14317 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n16559, B1 => 
                           REGISTERS_23_21_port, B2 => n16572, ZN => n16099);
   U14318 : NAND4_X1 port map( A1 => n16102, A2 => n16101, A3 => n16100, A4 => 
                           n16099, ZN => n16108);
   U14319 : AOI22_X1 port map( A1 => REGISTERS_19_21_port, A2 => n16569, B1 => 
                           REGISTERS_28_21_port, B2 => n16570, ZN => n16106);
   U14320 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n16557, B1 => 
                           REGISTERS_8_21_port, B2 => n16567, ZN => n16105);
   U14321 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n16574, B1 => 
                           REGISTERS_22_21_port, B2 => n16556, ZN => n16104);
   U14322 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n16580, B1 => 
                           REGISTERS_15_21_port, B2 => n16558, ZN => n16103);
   U14323 : NAND4_X1 port map( A1 => n16106, A2 => n16105, A3 => n16104, A4 => 
                           n16103, ZN => n16107);
   U14324 : NOR3_X1 port map( A1 => n16109, A2 => n16108, A3 => n16107, ZN => 
                           n16115);
   U14325 : AOI22_X1 port map( A1 => REGISTERS_2_21_port, A2 => n16545, B1 => 
                           REGISTERS_1_21_port, B2 => n16430, ZN => n16113);
   U14326 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n16542, B1 => 
                           REGISTERS_7_21_port, B2 => n16454, ZN => n16112);
   U14327 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n16597, B1 => 
                           REGISTERS_4_21_port, B2 => n16595, ZN => n16111);
   U14328 : AOI22_X1 port map( A1 => REGISTERS_3_21_port, A2 => n16593, B1 => 
                           REGISTERS_6_21_port, B2 => n16546, ZN => n16110);
   U14329 : OAI222_X1 port map( A1 => n15796, A2 => n16115, B1 => n16603, B2 =>
                           n16114, C1 => n14910, C2 => n8399, ZN => n8612);
   U14330 : AOI22_X1 port map( A1 => REGISTERS_23_20_port, A2 => n16572, B1 => 
                           REGISTERS_28_20_port, B2 => n16570, ZN => n16119);
   U14331 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n16557, B1 => 
                           REGISTERS_16_20_port, B2 => n16561, ZN => n16118);
   U14332 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n16567, B1 => 
                           REGISTERS_19_20_port, B2 => n16569, ZN => n16117);
   U14333 : AOI22_X1 port map( A1 => REGISTERS_30_20_port, A2 => n16555, B1 => 
                           REGISTERS_17_20_port, B2 => n16579, ZN => n16116);
   U14334 : NAND4_X1 port map( A1 => n16119, A2 => n16118, A3 => n16117, A4 => 
                           n16116, ZN => n16130);
   U14335 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n16574, B1 => 
                           REGISTERS_14_20_port, B2 => n16571, ZN => n16123);
   U14336 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n16562, B1 => 
                           REGISTERS_26_20_port, B2 => n16582, ZN => n16122);
   U14337 : AOI22_X1 port map( A1 => REGISTERS_18_20_port, A2 => n16584, B1 => 
                           REGISTERS_21_20_port, B2 => n16568, ZN => n16121);
   U14338 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n16581, B1 => 
                           REGISTERS_22_20_port, B2 => n16556, ZN => n16120);
   U14339 : NAND4_X1 port map( A1 => n16123, A2 => n16122, A3 => n16121, A4 => 
                           n16120, ZN => n16129);
   U14340 : AOI22_X1 port map( A1 => REGISTERS_27_20_port, A2 => n16573, B1 => 
                           REGISTERS_9_20_port, B2 => n16525, ZN => n16127);
   U14341 : AOI22_X1 port map( A1 => REGISTERS_10_20_port, A2 => n16560, B1 => 
                           REGISTERS_24_20_port, B2 => n16559, ZN => n16126);
   U14342 : AOI22_X1 port map( A1 => REGISTERS_31_20_port, A2 => n16583, B1 => 
                           REGISTERS_15_20_port, B2 => n16558, ZN => n16125);
   U14343 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n16580, B1 => 
                           REGISTERS_11_20_port, B2 => n15782, ZN => n16124);
   U14344 : NAND4_X1 port map( A1 => n16127, A2 => n16126, A3 => n16125, A4 => 
                           n16124, ZN => n16128);
   U14345 : NOR3_X1 port map( A1 => n16130, A2 => n16129, A3 => n16128, ZN => 
                           n16136);
   U14346 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n16595, B1 => 
                           REGISTERS_3_20_port, B2 => n16593, ZN => n16134);
   U14347 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n16542, B1 => 
                           REGISTERS_0_20_port, B2 => n16547, ZN => n16133);
   U14348 : AOI22_X1 port map( A1 => REGISTERS_2_20_port, A2 => n16545, B1 => 
                           REGISTERS_1_20_port, B2 => n16430, ZN => n16132);
   U14349 : AOI22_X1 port map( A1 => REGISTERS_7_20_port, A2 => n16454, B1 => 
                           REGISTERS_6_20_port, B2 => n16546, ZN => n16131);
   U14350 : AND4_X1 port map( A1 => n16134, A2 => n16133, A3 => n16132, A4 => 
                           n16131, ZN => n16135);
   U14351 : OAI222_X1 port map( A1 => n15796, A2 => n16136, B1 => n16603, B2 =>
                           n16135, C1 => n16071, C2 => n8398, ZN => n8613);
   U14352 : AOI22_X1 port map( A1 => REGISTERS_15_19_port, A2 => n16558, B1 => 
                           REGISTERS_24_19_port, B2 => n16559, ZN => n16140);
   U14353 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n16568, B1 => 
                           REGISTERS_28_19_port, B2 => n16570, ZN => n16139);
   U14354 : AOI22_X1 port map( A1 => REGISTERS_23_19_port, A2 => n16572, B1 => 
                           REGISTERS_8_19_port, B2 => n16567, ZN => n16138);
   U14355 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n16562, B1 => 
                           REGISTERS_18_19_port, B2 => n16584, ZN => n16137);
   U14356 : NAND4_X1 port map( A1 => n16140, A2 => n16139, A3 => n16138, A4 => 
                           n16137, ZN => n16151);
   U14357 : AOI22_X1 port map( A1 => REGISTERS_22_19_port, A2 => n16556, B1 => 
                           REGISTERS_20_19_port, B2 => n16581, ZN => n16144);
   U14358 : AOI22_X1 port map( A1 => REGISTERS_27_19_port, A2 => n16573, B1 => 
                           REGISTERS_12_19_port, B2 => n16580, ZN => n16143);
   U14359 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n16437, B1 => 
                           REGISTERS_25_19_port, B2 => n16557, ZN => n16142);
   U14360 : AOI22_X1 port map( A1 => REGISTERS_11_19_port, A2 => n15782, B1 => 
                           REGISTERS_31_19_port, B2 => n16583, ZN => n16141);
   U14361 : NAND4_X1 port map( A1 => n16144, A2 => n16143, A3 => n16142, A4 => 
                           n16141, ZN => n16150);
   U14362 : AOI22_X1 port map( A1 => REGISTERS_14_19_port, A2 => n16571, B1 => 
                           REGISTERS_30_19_port, B2 => n16555, ZN => n16148);
   U14363 : AOI22_X1 port map( A1 => REGISTERS_10_19_port, A2 => n16560, B1 => 
                           REGISTERS_26_19_port, B2 => n16582, ZN => n16147);
   U14364 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n16561, B1 => 
                           REGISTERS_19_19_port, B2 => n16569, ZN => n16146);
   U14365 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n16579, B1 => 
                           REGISTERS_29_19_port, B2 => n16574, ZN => n16145);
   U14366 : NAND4_X1 port map( A1 => n16148, A2 => n16147, A3 => n16146, A4 => 
                           n16145, ZN => n16149);
   U14367 : NOR3_X1 port map( A1 => n16151, A2 => n16150, A3 => n16149, ZN => 
                           n16157);
   U14368 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n16595, B1 => 
                           REGISTERS_6_19_port, B2 => n16546, ZN => n16155);
   U14369 : AOI22_X1 port map( A1 => REGISTERS_2_19_port, A2 => n16545, B1 => 
                           REGISTERS_0_19_port, B2 => n16547, ZN => n16154);
   U14370 : AOI22_X1 port map( A1 => REGISTERS_7_19_port, A2 => n16454, B1 => 
                           REGISTERS_3_19_port, B2 => n16593, ZN => n16153);
   U14371 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n16542, B1 => 
                           REGISTERS_1_19_port, B2 => n16430, ZN => n16152);
   U14372 : AND4_X1 port map( A1 => n16155, A2 => n16154, A3 => n16153, A4 => 
                           n16152, ZN => n16156);
   U14373 : OAI222_X1 port map( A1 => n16605, A2 => n16157, B1 => n16603, B2 =>
                           n16156, C1 => n14910, C2 => n8397, ZN => n8614);
   U14374 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n16562, B1 => 
                           REGISTERS_26_18_port, B2 => n16582, ZN => n16161);
   U14375 : AOI22_X1 port map( A1 => REGISTERS_23_18_port, A2 => n16572, B1 => 
                           REGISTERS_19_18_port, B2 => n16569, ZN => n16160);
   U14376 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n16581, B1 => 
                           REGISTERS_30_18_port, B2 => n16555, ZN => n16159);
   U14377 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n16559, B1 => 
                           REGISTERS_17_18_port, B2 => n16579, ZN => n16158);
   U14378 : NAND4_X1 port map( A1 => n16161, A2 => n16160, A3 => n16159, A4 => 
                           n16158, ZN => n16172);
   U14379 : AOI22_X1 port map( A1 => REGISTERS_31_18_port, A2 => n16583, B1 => 
                           REGISTERS_14_18_port, B2 => n16571, ZN => n16165);
   U14380 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n16561, B1 => 
                           REGISTERS_28_18_port, B2 => n16570, ZN => n16164);
   U14381 : AOI22_X1 port map( A1 => REGISTERS_27_18_port, A2 => n16573, B1 => 
                           REGISTERS_11_18_port, B2 => n16414, ZN => n16163);
   U14382 : AOI22_X1 port map( A1 => REGISTERS_18_18_port, A2 => n16584, B1 => 
                           REGISTERS_12_18_port, B2 => n16580, ZN => n16162);
   U14383 : NAND4_X1 port map( A1 => n16165, A2 => n16164, A3 => n16163, A4 => 
                           n16162, ZN => n16171);
   U14384 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n16567, B1 => 
                           REGISTERS_9_18_port, B2 => n16029, ZN => n16169);
   U14385 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n16568, B1 => 
                           REGISTERS_25_18_port, B2 => n16557, ZN => n16168);
   U14386 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n16574, B1 => 
                           REGISTERS_15_18_port, B2 => n16558, ZN => n16167);
   U14387 : AOI22_X1 port map( A1 => REGISTERS_10_18_port, A2 => n16560, B1 => 
                           REGISTERS_22_18_port, B2 => n16556, ZN => n16166);
   U14388 : NAND4_X1 port map( A1 => n16169, A2 => n16168, A3 => n16167, A4 => 
                           n16166, ZN => n16170);
   U14389 : NOR3_X1 port map( A1 => n16172, A2 => n16171, A3 => n16170, ZN => 
                           n16178);
   U14390 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n16597, B1 => 
                           REGISTERS_7_18_port, B2 => n16454, ZN => n16176);
   U14391 : AOI22_X1 port map( A1 => REGISTERS_6_18_port, A2 => n16344, B1 => 
                           REGISTERS_4_18_port, B2 => n16543, ZN => n16175);
   U14392 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n16544, B1 => 
                           REGISTERS_5_18_port, B2 => n16518, ZN => n16174);
   U14393 : AOI22_X1 port map( A1 => REGISTERS_2_18_port, A2 => n16545, B1 => 
                           REGISTERS_3_18_port, B2 => n16453, ZN => n16173);
   U14394 : AND4_X1 port map( A1 => n16176, A2 => n16175, A3 => n16174, A4 => 
                           n16173, ZN => n16177);
   U14395 : OAI222_X1 port map( A1 => n15796, A2 => n16178, B1 => n16603, B2 =>
                           n16177, C1 => n16071, C2 => n8396, ZN => n8615);
   U14396 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n16567, B1 => 
                           REGISTERS_13_17_port, B2 => n16562, ZN => n16182);
   U14397 : AOI22_X1 port map( A1 => REGISTERS_31_17_port, A2 => n16583, B1 => 
                           REGISTERS_30_17_port, B2 => n16555, ZN => n16181);
   U14398 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n16579, B1 => 
                           REGISTERS_19_17_port, B2 => n16569, ZN => n16180);
   U14399 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n16568, B1 => 
                           REGISTERS_11_17_port, B2 => n16414, ZN => n16179);
   U14400 : NAND4_X1 port map( A1 => n16182, A2 => n16181, A3 => n16180, A4 => 
                           n16179, ZN => n16193);
   U14401 : AOI22_X1 port map( A1 => REGISTERS_26_17_port, A2 => n16582, B1 => 
                           REGISTERS_18_17_port, B2 => n16584, ZN => n16186);
   U14402 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n16581, B1 => 
                           REGISTERS_27_17_port, B2 => n16573, ZN => n16185);
   U14403 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n16561, B1 => 
                           REGISTERS_14_17_port, B2 => n16571, ZN => n16184);
   U14404 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n16559, B1 => 
                           REGISTERS_9_17_port, B2 => n16525, ZN => n16183);
   U14405 : NAND4_X1 port map( A1 => n16186, A2 => n16185, A3 => n16184, A4 => 
                           n16183, ZN => n16192);
   U14406 : AOI22_X1 port map( A1 => REGISTERS_23_17_port, A2 => n16572, B1 => 
                           REGISTERS_29_17_port, B2 => n16574, ZN => n16190);
   U14407 : AOI22_X1 port map( A1 => REGISTERS_15_17_port, A2 => n16558, B1 => 
                           REGISTERS_10_17_port, B2 => n16560, ZN => n16189);
   U14408 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n16580, B1 => 
                           REGISTERS_28_17_port, B2 => n16570, ZN => n16188);
   U14409 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n16557, B1 => 
                           REGISTERS_22_17_port, B2 => n16556, ZN => n16187);
   U14410 : NAND4_X1 port map( A1 => n16190, A2 => n16189, A3 => n16188, A4 => 
                           n16187, ZN => n16191);
   U14411 : NOR3_X1 port map( A1 => n16193, A2 => n16192, A3 => n16191, ZN => 
                           n16199);
   U14412 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n16430, B1 => 
                           REGISTERS_5_17_port, B2 => n16518, ZN => n16197);
   U14413 : AOI22_X1 port map( A1 => REGISTERS_3_17_port, A2 => n16453, B1 => 
                           REGISTERS_6_17_port, B2 => n16546, ZN => n16196);
   U14414 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n16595, B1 => 
                           REGISTERS_2_17_port, B2 => n16596, ZN => n16195);
   U14415 : AOI22_X1 port map( A1 => REGISTERS_7_17_port, A2 => n16454, B1 => 
                           REGISTERS_0_17_port, B2 => n16547, ZN => n16194);
   U14416 : AND4_X1 port map( A1 => n16197, A2 => n16196, A3 => n16195, A4 => 
                           n16194, ZN => n16198);
   U14417 : OAI222_X1 port map( A1 => n16605, A2 => n16199, B1 => n16603, B2 =>
                           n16198, C1 => n16026, C2 => n8395, ZN => n8616);
   U14418 : AOI22_X1 port map( A1 => REGISTERS_15_16_port, A2 => n16558, B1 => 
                           REGISTERS_24_16_port, B2 => n16559, ZN => n16203);
   U14419 : AOI22_X1 port map( A1 => REGISTERS_18_16_port, A2 => n16584, B1 => 
                           REGISTERS_21_16_port, B2 => n16568, ZN => n16202);
   U14420 : AOI22_X1 port map( A1 => REGISTERS_30_16_port, A2 => n16555, B1 => 
                           REGISTERS_9_16_port, B2 => n16525, ZN => n16201);
   U14421 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n16581, B1 => 
                           REGISTERS_11_16_port, B2 => n16414, ZN => n16200);
   U14422 : NAND4_X1 port map( A1 => n16203, A2 => n16202, A3 => n16201, A4 => 
                           n16200, ZN => n16214);
   U14423 : AOI22_X1 port map( A1 => REGISTERS_31_16_port, A2 => n16583, B1 => 
                           REGISTERS_25_16_port, B2 => n16557, ZN => n16207);
   U14424 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n16567, B1 => 
                           REGISTERS_19_16_port, B2 => n16569, ZN => n16206);
   U14425 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n16580, B1 => 
                           REGISTERS_10_16_port, B2 => n16560, ZN => n16205);
   U14426 : AOI22_X1 port map( A1 => REGISTERS_14_16_port, A2 => n16571, B1 => 
                           REGISTERS_23_16_port, B2 => n16572, ZN => n16204);
   U14427 : NAND4_X1 port map( A1 => n16207, A2 => n16206, A3 => n16205, A4 => 
                           n16204, ZN => n16213);
   U14428 : AOI22_X1 port map( A1 => REGISTERS_22_16_port, A2 => n16556, B1 => 
                           REGISTERS_13_16_port, B2 => n16562, ZN => n16211);
   U14429 : AOI22_X1 port map( A1 => REGISTERS_26_16_port, A2 => n16582, B1 => 
                           REGISTERS_16_16_port, B2 => n16561, ZN => n16210);
   U14430 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n16579, B1 => 
                           REGISTERS_29_16_port, B2 => n16574, ZN => n16209);
   U14431 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n16570, B1 => 
                           REGISTERS_27_16_port, B2 => n16573, ZN => n16208);
   U14432 : NAND4_X1 port map( A1 => n16211, A2 => n16210, A3 => n16209, A4 => 
                           n16208, ZN => n16212);
   U14433 : NOR3_X1 port map( A1 => n16214, A2 => n16213, A3 => n16212, ZN => 
                           n16222);
   U14434 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n16322, B1 => 
                           REGISTERS_3_16_port, B2 => n16453, ZN => n16220);
   U14435 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n16597, B1 => 
                           REGISTERS_2_16_port, B2 => n16596, ZN => n16219);
   U14436 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n16215, B1 => 
                           REGISTERS_4_16_port, B2 => n16543, ZN => n16218);
   U14437 : AOI22_X1 port map( A1 => REGISTERS_7_16_port, A2 => n16216, B1 => 
                           REGISTERS_6_16_port, B2 => n16546, ZN => n16217);
   U14438 : AND4_X1 port map( A1 => n16220, A2 => n16219, A3 => n16218, A4 => 
                           n16217, ZN => n16221);
   U14439 : OAI222_X1 port map( A1 => n15796, A2 => n16222, B1 => n16603, B2 =>
                           n16221, C1 => n14910, C2 => n8394, ZN => n8617);
   U14440 : AOI22_X1 port map( A1 => REGISTERS_23_15_port, A2 => n16572, B1 => 
                           REGISTERS_16_15_port, B2 => n16561, ZN => n16226);
   U14441 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n16568, B1 => 
                           REGISTERS_11_15_port, B2 => n15782, ZN => n16225);
   U14442 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n16567, B1 => 
                           REGISTERS_19_15_port, B2 => n16569, ZN => n16224);
   U14443 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n16525, B1 => 
                           REGISTERS_13_15_port, B2 => n16562, ZN => n16223);
   U14444 : NAND4_X1 port map( A1 => n16226, A2 => n16225, A3 => n16224, A4 => 
                           n16223, ZN => n16237);
   U14445 : AOI22_X1 port map( A1 => REGISTERS_31_15_port, A2 => n16583, B1 => 
                           REGISTERS_12_15_port, B2 => n16580, ZN => n16230);
   U14446 : AOI22_X1 port map( A1 => REGISTERS_26_15_port, A2 => n16582, B1 => 
                           REGISTERS_24_15_port, B2 => n16559, ZN => n16229);
   U14447 : AOI22_X1 port map( A1 => REGISTERS_27_15_port, A2 => n16573, B1 => 
                           REGISTERS_30_15_port, B2 => n16555, ZN => n16228);
   U14448 : AOI22_X1 port map( A1 => REGISTERS_14_15_port, A2 => n16571, B1 => 
                           REGISTERS_25_15_port, B2 => n16557, ZN => n16227);
   U14449 : NAND4_X1 port map( A1 => n16230, A2 => n16229, A3 => n16228, A4 => 
                           n16227, ZN => n16236);
   U14450 : AOI22_X1 port map( A1 => REGISTERS_22_15_port, A2 => n16556, B1 => 
                           REGISTERS_18_15_port, B2 => n16584, ZN => n16234);
   U14451 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n16581, B1 => 
                           REGISTERS_15_15_port, B2 => n16558, ZN => n16233);
   U14452 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n16570, B1 => 
                           REGISTERS_10_15_port, B2 => n16560, ZN => n16232);
   U14453 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n16574, B1 => 
                           REGISTERS_17_15_port, B2 => n16579, ZN => n16231);
   U14454 : NAND4_X1 port map( A1 => n16234, A2 => n16233, A3 => n16232, A4 => 
                           n16231, ZN => n16235);
   U14455 : NOR3_X1 port map( A1 => n16237, A2 => n16236, A3 => n16235, ZN => 
                           n16243);
   U14456 : AOI22_X1 port map( A1 => REGISTERS_7_15_port, A2 => n16454, B1 => 
                           REGISTERS_5_15_port, B2 => n16518, ZN => n16241);
   U14457 : AOI22_X1 port map( A1 => REGISTERS_6_15_port, A2 => n16344, B1 => 
                           REGISTERS_0_15_port, B2 => n16547, ZN => n16240);
   U14458 : AOI22_X1 port map( A1 => REGISTERS_3_15_port, A2 => n16453, B1 => 
                           REGISTERS_2_15_port, B2 => n16596, ZN => n16239);
   U14459 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n16430, B1 => 
                           REGISTERS_4_15_port, B2 => n16543, ZN => n16238);
   U14460 : AND4_X1 port map( A1 => n16241, A2 => n16240, A3 => n16239, A4 => 
                           n16238, ZN => n16242);
   U14461 : OAI222_X1 port map( A1 => n16605, A2 => n16243, B1 => n16553, B2 =>
                           n16242, C1 => n16071, C2 => n8393, ZN => n8618);
   U14462 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n16561, B1 => 
                           REGISTERS_30_14_port, B2 => n16555, ZN => n16247);
   U14463 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n16525, B1 => 
                           REGISTERS_14_14_port, B2 => n16571, ZN => n16246);
   U14464 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n16580, B1 => 
                           REGISTERS_22_14_port, B2 => n16556, ZN => n16245);
   U14465 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n16581, B1 => 
                           REGISTERS_27_14_port, B2 => n16573, ZN => n16244);
   U14466 : NAND4_X1 port map( A1 => n16247, A2 => n16246, A3 => n16245, A4 => 
                           n16244, ZN => n16258);
   U14467 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n16568, B1 => 
                           REGISTERS_17_14_port, B2 => n16579, ZN => n16251);
   U14468 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n16559, B1 => 
                           REGISTERS_31_14_port, B2 => n16583, ZN => n16250);
   U14469 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n16562, B1 => 
                           REGISTERS_28_14_port, B2 => n16570, ZN => n16249);
   U14470 : AOI22_X1 port map( A1 => REGISTERS_26_14_port, A2 => n16582, B1 => 
                           REGISTERS_25_14_port, B2 => n16557, ZN => n16248);
   U14471 : NAND4_X1 port map( A1 => n16251, A2 => n16250, A3 => n16249, A4 => 
                           n16248, ZN => n16257);
   U14472 : AOI22_X1 port map( A1 => REGISTERS_19_14_port, A2 => n16569, B1 => 
                           REGISTERS_11_14_port, B2 => n16414, ZN => n16255);
   U14473 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n16574, B1 => 
                           REGISTERS_15_14_port, B2 => n16558, ZN => n16254);
   U14474 : AOI22_X1 port map( A1 => REGISTERS_10_14_port, A2 => n16560, B1 => 
                           REGISTERS_18_14_port, B2 => n16584, ZN => n16253);
   U14475 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n16567, B1 => 
                           REGISTERS_23_14_port, B2 => n16572, ZN => n16252);
   U14476 : NAND4_X1 port map( A1 => n16255, A2 => n16254, A3 => n16253, A4 => 
                           n16252, ZN => n16256);
   U14477 : NOR3_X1 port map( A1 => n16258, A2 => n16257, A3 => n16256, ZN => 
                           n16264);
   U14478 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n16595, B1 => 
                           REGISTERS_3_14_port, B2 => n16453, ZN => n16262);
   U14479 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n16322, B1 => 
                           REGISTERS_7_14_port, B2 => n16454, ZN => n16261);
   U14480 : AOI22_X1 port map( A1 => REGISTERS_2_14_port, A2 => n16545, B1 => 
                           REGISTERS_6_14_port, B2 => n16592, ZN => n16260);
   U14481 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n16542, B1 => 
                           REGISTERS_0_14_port, B2 => n16547, ZN => n16259);
   U14482 : AND4_X1 port map( A1 => n16262, A2 => n16261, A3 => n16260, A4 => 
                           n16259, ZN => n16263);
   U14483 : OAI222_X1 port map( A1 => n15796, A2 => n16264, B1 => n16553, B2 =>
                           n16263, C1 => n16026, C2 => n8392, ZN => n8619);
   U14484 : AOI22_X1 port map( A1 => REGISTERS_27_13_port, A2 => n16573, B1 => 
                           REGISTERS_30_13_port, B2 => n16555, ZN => n16268);
   U14485 : AOI22_X1 port map( A1 => REGISTERS_19_13_port, A2 => n16569, B1 => 
                           REGISTERS_13_13_port, B2 => n16562, ZN => n16267);
   U14486 : AOI22_X1 port map( A1 => REGISTERS_15_13_port, A2 => n16558, B1 => 
                           REGISTERS_14_13_port, B2 => n16571, ZN => n16266);
   U14487 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n16568, B1 => 
                           REGISTERS_25_13_port, B2 => n16557, ZN => n16265);
   U14488 : NAND4_X1 port map( A1 => n16268, A2 => n16267, A3 => n16266, A4 => 
                           n16265, ZN => n16279);
   U14489 : AOI22_X1 port map( A1 => REGISTERS_22_13_port, A2 => n16556, B1 => 
                           REGISTERS_31_13_port, B2 => n16583, ZN => n16272);
   U14490 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n16580, B1 => 
                           REGISTERS_8_13_port, B2 => n16567, ZN => n16271);
   U14491 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n16570, B1 => 
                           REGISTERS_29_13_port, B2 => n16574, ZN => n16270);
   U14492 : AOI22_X1 port map( A1 => REGISTERS_18_13_port, A2 => n16584, B1 => 
                           REGISTERS_16_13_port, B2 => n16561, ZN => n16269);
   U14493 : NAND4_X1 port map( A1 => n16272, A2 => n16271, A3 => n16270, A4 => 
                           n16269, ZN => n16278);
   U14494 : AOI22_X1 port map( A1 => REGISTERS_26_13_port, A2 => n16582, B1 => 
                           REGISTERS_9_13_port, B2 => n16029, ZN => n16276);
   U14495 : AOI22_X1 port map( A1 => REGISTERS_23_13_port, A2 => n16572, B1 => 
                           REGISTERS_20_13_port, B2 => n16581, ZN => n16275);
   U14496 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n16559, B1 => 
                           REGISTERS_10_13_port, B2 => n16560, ZN => n16274);
   U14497 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n16579, B1 => 
                           REGISTERS_11_13_port, B2 => n15782, ZN => n16273);
   U14498 : NAND4_X1 port map( A1 => n16276, A2 => n16275, A3 => n16274, A4 => 
                           n16273, ZN => n16277);
   U14499 : NOR3_X1 port map( A1 => n16279, A2 => n16278, A3 => n16277, ZN => 
                           n16285);
   U14500 : AOI22_X1 port map( A1 => REGISTERS_7_13_port, A2 => n16454, B1 => 
                           REGISTERS_5_13_port, B2 => n16518, ZN => n16283);
   U14501 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n16544, B1 => 
                           REGISTERS_2_13_port, B2 => n16596, ZN => n16282);
   U14502 : AOI22_X1 port map( A1 => REGISTERS_6_13_port, A2 => n16592, B1 => 
                           REGISTERS_3_13_port, B2 => n16453, ZN => n16281);
   U14503 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n16597, B1 => 
                           REGISTERS_4_13_port, B2 => n16543, ZN => n16280);
   U14504 : OAI222_X1 port map( A1 => n16605, A2 => n16285, B1 => n16603, B2 =>
                           n16284, C1 => n14910, C2 => n8391, ZN => n8620);
   U14505 : AOI22_X1 port map( A1 => REGISTERS_27_12_port, A2 => n16573, B1 => 
                           REGISTERS_26_12_port, B2 => n16582, ZN => n16289);
   U14506 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n16568, B1 => 
                           REGISTERS_20_12_port, B2 => n16581, ZN => n16288);
   U14507 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n16559, B1 => 
                           REGISTERS_25_12_port, B2 => n16557, ZN => n16287);
   U14508 : AOI22_X1 port map( A1 => REGISTERS_23_12_port, A2 => n16572, B1 => 
                           REGISTERS_19_12_port, B2 => n16569, ZN => n16286);
   U14509 : NAND4_X1 port map( A1 => n16289, A2 => n16288, A3 => n16287, A4 => 
                           n16286, ZN => n16300);
   U14510 : AOI22_X1 port map( A1 => REGISTERS_11_12_port, A2 => n16530, B1 => 
                           REGISTERS_29_12_port, B2 => n16574, ZN => n16293);
   U14511 : AOI22_X1 port map( A1 => REGISTERS_10_12_port, A2 => n16560, B1 => 
                           REGISTERS_16_12_port, B2 => n16561, ZN => n16292);
   U14512 : AOI22_X1 port map( A1 => REGISTERS_18_12_port, A2 => n16584, B1 => 
                           REGISTERS_9_12_port, B2 => n16525, ZN => n16291);
   U14513 : AOI22_X1 port map( A1 => REGISTERS_15_12_port, A2 => n16558, B1 => 
                           REGISTERS_13_12_port, B2 => n16562, ZN => n16290);
   U14514 : NAND4_X1 port map( A1 => n16293, A2 => n16292, A3 => n16291, A4 => 
                           n16290, ZN => n16299);
   U14515 : AOI22_X1 port map( A1 => REGISTERS_31_12_port, A2 => n16583, B1 => 
                           REGISTERS_30_12_port, B2 => n16555, ZN => n16297);
   U14516 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n16567, B1 => 
                           REGISTERS_28_12_port, B2 => n16570, ZN => n16296);
   U14517 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n16580, B1 => 
                           REGISTERS_17_12_port, B2 => n16579, ZN => n16295);
   U14518 : AOI22_X1 port map( A1 => REGISTERS_14_12_port, A2 => n16571, B1 => 
                           REGISTERS_22_12_port, B2 => n16556, ZN => n16294);
   U14519 : NAND4_X1 port map( A1 => n16297, A2 => n16296, A3 => n16295, A4 => 
                           n16294, ZN => n16298);
   U14520 : NOR3_X1 port map( A1 => n16300, A2 => n16299, A3 => n16298, ZN => 
                           n16306);
   U14521 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n16595, B1 => 
                           REGISTERS_7_12_port, B2 => n16454, ZN => n16304);
   U14522 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n16544, B1 => 
                           REGISTERS_2_12_port, B2 => n16596, ZN => n16303);
   U14523 : AOI22_X1 port map( A1 => REGISTERS_3_12_port, A2 => n16593, B1 => 
                           REGISTERS_5_12_port, B2 => n16518, ZN => n16302);
   U14524 : AOI22_X1 port map( A1 => REGISTERS_0_12_port, A2 => n16597, B1 => 
                           REGISTERS_6_12_port, B2 => n16592, ZN => n16301);
   U14525 : AND4_X1 port map( A1 => n16304, A2 => n16303, A3 => n16302, A4 => 
                           n16301, ZN => n16305);
   U14526 : OAI222_X1 port map( A1 => n15796, A2 => n16306, B1 => n16603, B2 =>
                           n16305, C1 => n16049, C2 => n8390, ZN => n8621);
   U14527 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n16568, B1 => 
                           REGISTERS_15_11_port, B2 => n16558, ZN => n16310);
   U14528 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n16561, B1 => 
                           REGISTERS_27_11_port, B2 => n16573, ZN => n16309);
   U14529 : AOI22_X1 port map( A1 => REGISTERS_23_11_port, A2 => n16572, B1 => 
                           REGISTERS_22_11_port, B2 => n16556, ZN => n16308);
   U14530 : AOI22_X1 port map( A1 => REGISTERS_10_11_port, A2 => n16560, B1 => 
                           REGISTERS_29_11_port, B2 => n16574, ZN => n16307);
   U14531 : NAND4_X1 port map( A1 => n16310, A2 => n16309, A3 => n16308, A4 => 
                           n16307, ZN => n16321);
   U14532 : AOI22_X1 port map( A1 => REGISTERS_31_11_port, A2 => n16583, B1 => 
                           REGISTERS_11_11_port, B2 => n16414, ZN => n16314);
   U14533 : AOI22_X1 port map( A1 => REGISTERS_14_11_port, A2 => n16571, B1 => 
                           REGISTERS_24_11_port, B2 => n16559, ZN => n16313);
   U14534 : AOI22_X1 port map( A1 => REGISTERS_18_11_port, A2 => n16584, B1 => 
                           REGISTERS_28_11_port, B2 => n16570, ZN => n16312);
   U14535 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n16567, B1 => 
                           REGISTERS_9_11_port, B2 => n16525, ZN => n16311);
   U14536 : NAND4_X1 port map( A1 => n16314, A2 => n16313, A3 => n16312, A4 => 
                           n16311, ZN => n16320);
   U14537 : AOI22_X1 port map( A1 => REGISTERS_19_11_port, A2 => n16569, B1 => 
                           REGISTERS_12_11_port, B2 => n16580, ZN => n16318);
   U14538 : AOI22_X1 port map( A1 => REGISTERS_26_11_port, A2 => n16582, B1 => 
                           REGISTERS_30_11_port, B2 => n16555, ZN => n16317);
   U14539 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n16579, B1 => 
                           REGISTERS_25_11_port, B2 => n16557, ZN => n16316);
   U14540 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n16581, B1 => 
                           REGISTERS_13_11_port, B2 => n16562, ZN => n16315);
   U14541 : NAND4_X1 port map( A1 => n16318, A2 => n16317, A3 => n16316, A4 => 
                           n16315, ZN => n16319);
   U14542 : NOR3_X1 port map( A1 => n16321, A2 => n16320, A3 => n16319, ZN => 
                           n16328);
   U14543 : AOI22_X1 port map( A1 => REGISTERS_2_11_port, A2 => n16545, B1 => 
                           REGISTERS_7_11_port, B2 => n16454, ZN => n16326);
   U14544 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n16322, B1 => 
                           REGISTERS_5_11_port, B2 => n16518, ZN => n16325);
   U14545 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n16597, B1 => 
                           REGISTERS_6_11_port, B2 => n16592, ZN => n16324);
   U14546 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n16595, B1 => 
                           REGISTERS_3_11_port, B2 => n16453, ZN => n16323);
   U14547 : AND4_X1 port map( A1 => n16326, A2 => n16325, A3 => n16324, A4 => 
                           n16323, ZN => n16327);
   U14548 : OAI222_X1 port map( A1 => n15796, A2 => n16328, B1 => n16553, B2 =>
                           n16327, C1 => n16071, C2 => n8389, ZN => n8622);
   U14549 : AOI22_X1 port map( A1 => REGISTERS_22_10_port, A2 => n16556, B1 => 
                           REGISTERS_16_10_port, B2 => n16561, ZN => n16332);
   U14550 : AOI22_X1 port map( A1 => REGISTERS_31_10_port, A2 => n16583, B1 => 
                           REGISTERS_8_10_port, B2 => n16567, ZN => n16331);
   U14551 : AOI22_X1 port map( A1 => REGISTERS_11_10_port, A2 => n16414, B1 => 
                           REGISTERS_15_10_port, B2 => n16558, ZN => n16330);
   U14552 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n16557, B1 => 
                           REGISTERS_19_10_port, B2 => n16569, ZN => n16329);
   U14553 : NAND4_X1 port map( A1 => n16332, A2 => n16331, A3 => n16330, A4 => 
                           n16329, ZN => n16343);
   U14554 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n16574, B1 => 
                           REGISTERS_20_10_port, B2 => n16581, ZN => n16336);
   U14555 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n16579, B1 => 
                           REGISTERS_13_10_port, B2 => n16562, ZN => n16335);
   U14556 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n16568, B1 => 
                           REGISTERS_28_10_port, B2 => n16570, ZN => n16334);
   U14557 : AOI22_X1 port map( A1 => REGISTERS_27_10_port, A2 => n16573, B1 => 
                           REGISTERS_30_10_port, B2 => n16555, ZN => n16333);
   U14558 : NAND4_X1 port map( A1 => n16336, A2 => n16335, A3 => n16334, A4 => 
                           n16333, ZN => n16342);
   U14559 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n16580, B1 => 
                           REGISTERS_9_10_port, B2 => n16525, ZN => n16340);
   U14560 : AOI22_X1 port map( A1 => REGISTERS_23_10_port, A2 => n16572, B1 => 
                           REGISTERS_26_10_port, B2 => n16582, ZN => n16339);
   U14561 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n16559, B1 => 
                           REGISTERS_18_10_port, B2 => n16584, ZN => n16338);
   U14562 : AOI22_X1 port map( A1 => REGISTERS_14_10_port, A2 => n16571, B1 => 
                           REGISTERS_10_10_port, B2 => n16560, ZN => n16337);
   U14563 : NAND4_X1 port map( A1 => n16340, A2 => n16339, A3 => n16338, A4 => 
                           n16337, ZN => n16341);
   U14564 : NOR3_X1 port map( A1 => n16343, A2 => n16342, A3 => n16341, ZN => 
                           n16350);
   U14565 : AOI22_X1 port map( A1 => REGISTERS_7_10_port, A2 => n16454, B1 => 
                           REGISTERS_0_10_port, B2 => n16547, ZN => n16348);
   U14566 : AOI22_X1 port map( A1 => REGISTERS_6_10_port, A2 => n16344, B1 => 
                           REGISTERS_2_10_port, B2 => n16596, ZN => n16347);
   U14567 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n16542, B1 => 
                           REGISTERS_1_10_port, B2 => n16544, ZN => n16346);
   U14568 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n16595, B1 => 
                           REGISTERS_3_10_port, B2 => n16453, ZN => n16345);
   U14569 : AND4_X1 port map( A1 => n16348, A2 => n16347, A3 => n16346, A4 => 
                           n16345, ZN => n16349);
   U14570 : OAI222_X1 port map( A1 => n16605, A2 => n16350, B1 => n16603, B2 =>
                           n16349, C1 => n16071, C2 => n8388, ZN => n8623);
   U14571 : AOI22_X1 port map( A1 => REGISTERS_23_9_port, A2 => n16572, B1 => 
                           REGISTERS_9_9_port, B2 => n16525, ZN => n16354);
   U14572 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n16562, B1 => 
                           REGISTERS_8_9_port, B2 => n16567, ZN => n16353);
   U14573 : AOI22_X1 port map( A1 => REGISTERS_26_9_port, A2 => n16582, B1 => 
                           REGISTERS_24_9_port, B2 => n16559, ZN => n16352);
   U14574 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n16581, B1 => 
                           REGISTERS_15_9_port, B2 => n16558, ZN => n16351);
   U14575 : NAND4_X1 port map( A1 => n16354, A2 => n16353, A3 => n16352, A4 => 
                           n16351, ZN => n16365);
   U14576 : AOI22_X1 port map( A1 => REGISTERS_31_9_port, A2 => n16583, B1 => 
                           REGISTERS_30_9_port, B2 => n16555, ZN => n16358);
   U14577 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n16580, B1 => 
                           REGISTERS_17_9_port, B2 => n16579, ZN => n16357);
   U14578 : AOI22_X1 port map( A1 => REGISTERS_11_9_port, A2 => n16414, B1 => 
                           REGISTERS_14_9_port, B2 => n16571, ZN => n16356);
   U14579 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n16570, B1 => 
                           REGISTERS_25_9_port, B2 => n16557, ZN => n16355);
   U14580 : NAND4_X1 port map( A1 => n16358, A2 => n16357, A3 => n16356, A4 => 
                           n16355, ZN => n16364);
   U14581 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n16568, B1 => 
                           REGISTERS_19_9_port, B2 => n16569, ZN => n16362);
   U14582 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n16561, B1 => 
                           REGISTERS_22_9_port, B2 => n16556, ZN => n16361);
   U14583 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n16574, B1 => 
                           REGISTERS_27_9_port, B2 => n16573, ZN => n16360);
   U14584 : AOI22_X1 port map( A1 => REGISTERS_18_9_port, A2 => n16584, B1 => 
                           REGISTERS_10_9_port, B2 => n16560, ZN => n16359);
   U14585 : NAND4_X1 port map( A1 => n16362, A2 => n16361, A3 => n16360, A4 => 
                           n16359, ZN => n16363);
   U14586 : NOR3_X1 port map( A1 => n16365, A2 => n16364, A3 => n16363, ZN => 
                           n16371);
   U14587 : AOI22_X1 port map( A1 => REGISTERS_7_9_port, A2 => n16454, B1 => 
                           REGISTERS_1_9_port, B2 => n16544, ZN => n16369);
   U14588 : AOI22_X1 port map( A1 => REGISTERS_2_9_port, A2 => n16545, B1 => 
                           REGISTERS_0_9_port, B2 => n16547, ZN => n16368);
   U14589 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n16542, B1 => 
                           REGISTERS_6_9_port, B2 => n16592, ZN => n16367);
   U14590 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n16595, B1 => 
                           REGISTERS_3_9_port, B2 => n16453, ZN => n16366);
   U14591 : AND4_X1 port map( A1 => n16369, A2 => n16368, A3 => n16367, A4 => 
                           n16366, ZN => n16370);
   U14592 : OAI222_X1 port map( A1 => n15796, A2 => n16371, B1 => n16553, B2 =>
                           n16370, C1 => n16026, C2 => n8387, ZN => n8624);
   U14593 : AOI22_X1 port map( A1 => REGISTERS_10_8_port, A2 => n16560, B1 => 
                           REGISTERS_23_8_port, B2 => n16572, ZN => n16375);
   U14594 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n16437, B1 => 
                           REGISTERS_13_8_port, B2 => n16562, ZN => n16374);
   U14595 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n16579, B1 => 
                           REGISTERS_14_8_port, B2 => n16571, ZN => n16373);
   U14596 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n16561, B1 => 
                           REGISTERS_25_8_port, B2 => n16557, ZN => n16372);
   U14597 : NAND4_X1 port map( A1 => n16375, A2 => n16374, A3 => n16373, A4 => 
                           n16372, ZN => n16386);
   U14598 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n16574, B1 => 
                           REGISTERS_21_8_port, B2 => n16568, ZN => n16379);
   U14599 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n16570, B1 => 
                           REGISTERS_20_8_port, B2 => n16581, ZN => n16378);
   U14600 : AOI22_X1 port map( A1 => REGISTERS_26_8_port, A2 => n16582, B1 => 
                           REGISTERS_22_8_port, B2 => n16556, ZN => n16377);
   U14601 : AOI22_X1 port map( A1 => REGISTERS_31_8_port, A2 => n16583, B1 => 
                           REGISTERS_12_8_port, B2 => n16580, ZN => n16376);
   U14602 : NAND4_X1 port map( A1 => n16379, A2 => n16378, A3 => n16377, A4 => 
                           n16376, ZN => n16385);
   U14603 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n16559, B1 => 
                           REGISTERS_30_8_port, B2 => n16555, ZN => n16383);
   U14604 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n16567, B1 => 
                           REGISTERS_19_8_port, B2 => n16569, ZN => n16382);
   U14605 : AOI22_X1 port map( A1 => REGISTERS_27_8_port, A2 => n16573, B1 => 
                           REGISTERS_18_8_port, B2 => n16584, ZN => n16381);
   U14606 : AOI22_X1 port map( A1 => REGISTERS_11_8_port, A2 => n16414, B1 => 
                           REGISTERS_15_8_port, B2 => n16558, ZN => n16380);
   U14607 : NAND4_X1 port map( A1 => n16383, A2 => n16382, A3 => n16381, A4 => 
                           n16380, ZN => n16384);
   U14608 : NOR3_X1 port map( A1 => n16386, A2 => n16385, A3 => n16384, ZN => 
                           n16392);
   U14609 : AOI22_X1 port map( A1 => REGISTERS_2_8_port, A2 => n16545, B1 => 
                           REGISTERS_3_8_port, B2 => n16453, ZN => n16390);
   U14610 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n16595, B1 => 
                           REGISTERS_0_8_port, B2 => n16547, ZN => n16389);
   U14611 : AOI22_X1 port map( A1 => REGISTERS_7_8_port, A2 => n16454, B1 => 
                           REGISTERS_6_8_port, B2 => n16592, ZN => n16388);
   U14612 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n16542, B1 => 
                           REGISTERS_1_8_port, B2 => n16544, ZN => n16387);
   U14613 : AND4_X1 port map( A1 => n16390, A2 => n16389, A3 => n16388, A4 => 
                           n16387, ZN => n16391);
   U14614 : OAI222_X1 port map( A1 => n16605, A2 => n16392, B1 => n16603, B2 =>
                           n16391, C1 => n14910, C2 => n8386, ZN => n8625);
   U14615 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n16579, B1 => 
                           REGISTERS_14_7_port, B2 => n16571, ZN => n16396);
   U14616 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n16559, B1 => 
                           REGISTERS_25_7_port, B2 => n16557, ZN => n16395);
   U14617 : AOI22_X1 port map( A1 => REGISTERS_27_7_port, A2 => n16573, B1 => 
                           REGISTERS_30_7_port, B2 => n16555, ZN => n16394);
   U14618 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n16581, B1 => 
                           REGISTERS_8_7_port, B2 => n16567, ZN => n16393);
   U14619 : NAND4_X1 port map( A1 => n16396, A2 => n16395, A3 => n16394, A4 => 
                           n16393, ZN => n16407);
   U14620 : AOI22_X1 port map( A1 => REGISTERS_11_7_port, A2 => n16530, B1 => 
                           REGISTERS_23_7_port, B2 => n16572, ZN => n16400);
   U14621 : AOI22_X1 port map( A1 => REGISTERS_18_7_port, A2 => n16584, B1 => 
                           REGISTERS_26_7_port, B2 => n16582, ZN => n16399);
   U14622 : AOI22_X1 port map( A1 => REGISTERS_22_7_port, A2 => n16556, B1 => 
                           REGISTERS_9_7_port, B2 => n16525, ZN => n16398);
   U14623 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n16568, B1 => 
                           REGISTERS_16_7_port, B2 => n16561, ZN => n16397);
   U14624 : NAND4_X1 port map( A1 => n16400, A2 => n16399, A3 => n16398, A4 => 
                           n16397, ZN => n16406);
   U14625 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n16580, B1 => 
                           REGISTERS_28_7_port, B2 => n16570, ZN => n16404);
   U14626 : AOI22_X1 port map( A1 => REGISTERS_10_7_port, A2 => n16560, B1 => 
                           REGISTERS_15_7_port, B2 => n16558, ZN => n16403);
   U14627 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n16562, B1 => 
                           REGISTERS_19_7_port, B2 => n16569, ZN => n16402);
   U14628 : AOI22_X1 port map( A1 => REGISTERS_31_7_port, A2 => n16583, B1 => 
                           REGISTERS_29_7_port, B2 => n16574, ZN => n16401);
   U14629 : NAND4_X1 port map( A1 => n16404, A2 => n16403, A3 => n16402, A4 => 
                           n16401, ZN => n16405);
   U14630 : NOR3_X1 port map( A1 => n16407, A2 => n16406, A3 => n16405, ZN => 
                           n16413);
   U14631 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n16597, B1 => 
                           REGISTERS_5_7_port, B2 => n16518, ZN => n16411);
   U14632 : AOI22_X1 port map( A1 => REGISTERS_6_7_port, A2 => n16546, B1 => 
                           REGISTERS_1_7_port, B2 => n16430, ZN => n16410);
   U14633 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n16595, B1 => 
                           REGISTERS_3_7_port, B2 => n16453, ZN => n16409);
   U14634 : AOI22_X1 port map( A1 => REGISTERS_7_7_port, A2 => n16454, B1 => 
                           REGISTERS_2_7_port, B2 => n16596, ZN => n16408);
   U14635 : AND4_X1 port map( A1 => n16411, A2 => n16410, A3 => n16409, A4 => 
                           n16408, ZN => n16412);
   U14636 : OAI222_X1 port map( A1 => n15796, A2 => n16413, B1 => n16553, B2 =>
                           n16412, C1 => n16049, C2 => n8385, ZN => n8626);
   U14637 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n16568, B1 => 
                           REGISTERS_19_6_port, B2 => n16569, ZN => n16418);
   U14638 : AOI22_X1 port map( A1 => REGISTERS_15_6_port, A2 => n16558, B1 => 
                           REGISTERS_9_6_port, B2 => n16525, ZN => n16417);
   U14639 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n16567, B1 => 
                           REGISTERS_30_6_port, B2 => n16555, ZN => n16416);
   U14640 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n16580, B1 => 
                           REGISTERS_11_6_port, B2 => n16414, ZN => n16415);
   U14641 : NAND4_X1 port map( A1 => n16418, A2 => n16417, A3 => n16416, A4 => 
                           n16415, ZN => n16429);
   U14642 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n16581, B1 => 
                           REGISTERS_24_6_port, B2 => n16559, ZN => n16422);
   U14643 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n16557, B1 => 
                           REGISTERS_22_6_port, B2 => n16556, ZN => n16421);
   U14644 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n16579, B1 => 
                           REGISTERS_26_6_port, B2 => n16582, ZN => n16420);
   U14645 : AOI22_X1 port map( A1 => REGISTERS_10_6_port, A2 => n16560, B1 => 
                           REGISTERS_16_6_port, B2 => n16561, ZN => n16419);
   U14646 : NAND4_X1 port map( A1 => n16422, A2 => n16421, A3 => n16420, A4 => 
                           n16419, ZN => n16428);
   U14647 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n16570, B1 => 
                           REGISTERS_13_6_port, B2 => n16562, ZN => n16426);
   U14648 : AOI22_X1 port map( A1 => REGISTERS_23_6_port, A2 => n16572, B1 => 
                           REGISTERS_31_6_port, B2 => n16583, ZN => n16425);
   U14649 : AOI22_X1 port map( A1 => REGISTERS_14_6_port, A2 => n16571, B1 => 
                           REGISTERS_18_6_port, B2 => n16584, ZN => n16424);
   U14650 : AOI22_X1 port map( A1 => REGISTERS_27_6_port, A2 => n16573, B1 => 
                           REGISTERS_29_6_port, B2 => n16574, ZN => n16423);
   U14651 : NAND4_X1 port map( A1 => n16426, A2 => n16425, A3 => n16424, A4 => 
                           n16423, ZN => n16427);
   U14652 : NOR3_X1 port map( A1 => n16429, A2 => n16428, A3 => n16427, ZN => 
                           n16436);
   U14653 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n16595, B1 => 
                           REGISTERS_3_6_port, B2 => n16453, ZN => n16434);
   U14654 : AOI22_X1 port map( A1 => REGISTERS_6_6_port, A2 => n16546, B1 => 
                           REGISTERS_0_6_port, B2 => n16547, ZN => n16433);
   U14655 : AOI22_X1 port map( A1 => REGISTERS_2_6_port, A2 => n16545, B1 => 
                           REGISTERS_5_6_port, B2 => n16518, ZN => n16432);
   U14656 : AOI22_X1 port map( A1 => REGISTERS_7_6_port, A2 => n16454, B1 => 
                           REGISTERS_1_6_port, B2 => n16430, ZN => n16431);
   U14657 : OAI222_X1 port map( A1 => n16605, A2 => n16436, B1 => n16603, B2 =>
                           n16435, C1 => n16026, C2 => n8384, ZN => n8627);
   U14658 : AOI22_X1 port map( A1 => REGISTERS_15_5_port, A2 => n16558, B1 => 
                           REGISTERS_26_5_port, B2 => n16582, ZN => n16441);
   U14659 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n16557, B1 => 
                           REGISTERS_16_5_port, B2 => n16561, ZN => n16440);
   U14660 : AOI22_X1 port map( A1 => REGISTERS_11_5_port, A2 => n16530, B1 => 
                           REGISTERS_31_5_port, B2 => n16583, ZN => n16439);
   U14661 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n16437, B1 => 
                           REGISTERS_14_5_port, B2 => n16571, ZN => n16438);
   U14662 : NAND4_X1 port map( A1 => n16441, A2 => n16440, A3 => n16439, A4 => 
                           n16438, ZN => n16452);
   U14663 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n16568, B1 => 
                           REGISTERS_23_5_port, B2 => n16572, ZN => n16445);
   U14664 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n16567, B1 => 
                           REGISTERS_20_5_port, B2 => n16581, ZN => n16444);
   U14665 : AOI22_X1 port map( A1 => REGISTERS_10_5_port, A2 => n16560, B1 => 
                           REGISTERS_27_5_port, B2 => n16573, ZN => n16443);
   U14666 : AOI22_X1 port map( A1 => REGISTERS_30_5_port, A2 => n16555, B1 => 
                           REGISTERS_29_5_port, B2 => n16574, ZN => n16442);
   U14667 : NAND4_X1 port map( A1 => n16445, A2 => n16444, A3 => n16443, A4 => 
                           n16442, ZN => n16451);
   U14668 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n16562, B1 => 
                           REGISTERS_24_5_port, B2 => n16559, ZN => n16449);
   U14669 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n16570, B1 => 
                           REGISTERS_17_5_port, B2 => n16579, ZN => n16448);
   U14670 : AOI22_X1 port map( A1 => REGISTERS_22_5_port, A2 => n16556, B1 => 
                           REGISTERS_12_5_port, B2 => n16580, ZN => n16447);
   U14671 : AOI22_X1 port map( A1 => REGISTERS_19_5_port, A2 => n16569, B1 => 
                           REGISTERS_18_5_port, B2 => n16584, ZN => n16446);
   U14672 : NAND4_X1 port map( A1 => n16449, A2 => n16448, A3 => n16447, A4 => 
                           n16446, ZN => n16450);
   U14673 : NOR3_X1 port map( A1 => n16452, A2 => n16451, A3 => n16450, ZN => 
                           n16460);
   U14674 : AOI22_X1 port map( A1 => REGISTERS_0_5_port, A2 => n16597, B1 => 
                           REGISTERS_5_5_port, B2 => n16518, ZN => n16458);
   U14675 : AOI22_X1 port map( A1 => REGISTERS_3_5_port, A2 => n16453, B1 => 
                           REGISTERS_6_5_port, B2 => n16546, ZN => n16457);
   U14676 : AOI22_X1 port map( A1 => REGISTERS_7_5_port, A2 => n16454, B1 => 
                           REGISTERS_2_5_port, B2 => n16596, ZN => n16456);
   U14677 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n16544, B1 => 
                           REGISTERS_4_5_port, B2 => n16543, ZN => n16455);
   U14678 : AND4_X1 port map( A1 => n16458, A2 => n16457, A3 => n16456, A4 => 
                           n16455, ZN => n16459);
   U14679 : OAI222_X1 port map( A1 => n15796, A2 => n16460, B1 => n16553, B2 =>
                           n16459, C1 => n16071, C2 => n8383, ZN => n8628);
   U14680 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n16561, B1 => 
                           REGISTERS_29_4_port, B2 => n16574, ZN => n16464);
   U14681 : AOI22_X1 port map( A1 => REGISTERS_31_4_port, A2 => n16583, B1 => 
                           REGISTERS_27_4_port, B2 => n16573, ZN => n16463);
   U14682 : AOI22_X1 port map( A1 => REGISTERS_14_4_port, A2 => n16571, B1 => 
                           REGISTERS_21_4_port, B2 => n16568, ZN => n16462);
   U14683 : AOI22_X1 port map( A1 => REGISTERS_30_4_port, A2 => n16555, B1 => 
                           REGISTERS_24_4_port, B2 => n16559, ZN => n16461);
   U14684 : NAND4_X1 port map( A1 => n16464, A2 => n16463, A3 => n16462, A4 => 
                           n16461, ZN => n16475);
   U14685 : AOI22_X1 port map( A1 => REGISTERS_15_4_port, A2 => n16558, B1 => 
                           REGISTERS_10_4_port, B2 => n16560, ZN => n16468);
   U14686 : AOI22_X1 port map( A1 => REGISTERS_26_4_port, A2 => n16582, B1 => 
                           REGISTERS_22_4_port, B2 => n16556, ZN => n16467);
   U14687 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n16570, B1 => 
                           REGISTERS_19_4_port, B2 => n16569, ZN => n16466);
   U14688 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n16581, B1 => 
                           REGISTERS_23_4_port, B2 => n16572, ZN => n16465);
   U14689 : NAND4_X1 port map( A1 => n16468, A2 => n16467, A3 => n16466, A4 => 
                           n16465, ZN => n16474);
   U14690 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n16579, B1 => 
                           REGISTERS_18_4_port, B2 => n16584, ZN => n16472);
   U14691 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n16029, B1 => 
                           REGISTERS_12_4_port, B2 => n16580, ZN => n16471);
   U14692 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n16557, B1 => 
                           REGISTERS_8_4_port, B2 => n16567, ZN => n16470);
   U14693 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n16562, B1 => 
                           REGISTERS_11_4_port, B2 => n15782, ZN => n16469);
   U14694 : NAND4_X1 port map( A1 => n16472, A2 => n16471, A3 => n16470, A4 => 
                           n16469, ZN => n16473);
   U14695 : NOR3_X1 port map( A1 => n16475, A2 => n16474, A3 => n16473, ZN => 
                           n16481);
   U14696 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n16542, B1 => 
                           REGISTERS_7_4_port, B2 => n16454, ZN => n16479);
   U14697 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n16544, B1 => 
                           REGISTERS_3_4_port, B2 => n16593, ZN => n16478);
   U14698 : AOI22_X1 port map( A1 => REGISTERS_0_4_port, A2 => n16597, B1 => 
                           REGISTERS_4_4_port, B2 => n16543, ZN => n16477);
   U14699 : AOI22_X1 port map( A1 => REGISTERS_2_4_port, A2 => n16545, B1 => 
                           REGISTERS_6_4_port, B2 => n16546, ZN => n16476);
   U14700 : AND4_X1 port map( A1 => n16479, A2 => n16478, A3 => n16477, A4 => 
                           n16476, ZN => n16480);
   U14701 : OAI222_X1 port map( A1 => n16605, A2 => n16481, B1 => n16603, B2 =>
                           n16480, C1 => n16026, C2 => n8382, ZN => n8629);
   U14702 : AOI22_X1 port map( A1 => REGISTERS_14_3_port, A2 => n16571, B1 => 
                           REGISTERS_23_3_port, B2 => n16572, ZN => n16485);
   U14703 : AOI22_X1 port map( A1 => REGISTERS_31_3_port, A2 => n16583, B1 => 
                           REGISTERS_20_3_port, B2 => n16581, ZN => n16484);
   U14704 : AOI22_X1 port map( A1 => REGISTERS_22_3_port, A2 => n16556, B1 => 
                           REGISTERS_12_3_port, B2 => n16580, ZN => n16483);
   U14705 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n16567, B1 => 
                           REGISTERS_9_3_port, B2 => n16525, ZN => n16482);
   U14706 : NAND4_X1 port map( A1 => n16485, A2 => n16484, A3 => n16483, A4 => 
                           n16482, ZN => n16496);
   U14707 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n16559, B1 => 
                           REGISTERS_11_3_port, B2 => n16414, ZN => n16489);
   U14708 : AOI22_X1 port map( A1 => REGISTERS_30_3_port, A2 => n16555, B1 => 
                           REGISTERS_15_3_port, B2 => n16558, ZN => n16488);
   U14709 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n16562, B1 => 
                           REGISTERS_16_3_port, B2 => n16561, ZN => n16487);
   U14710 : AOI22_X1 port map( A1 => REGISTERS_27_3_port, A2 => n16573, B1 => 
                           REGISTERS_29_3_port, B2 => n16574, ZN => n16486);
   U14711 : NAND4_X1 port map( A1 => n16489, A2 => n16488, A3 => n16487, A4 => 
                           n16486, ZN => n16495);
   U14712 : AOI22_X1 port map( A1 => REGISTERS_26_3_port, A2 => n16582, B1 => 
                           REGISTERS_28_3_port, B2 => n16570, ZN => n16493);
   U14713 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n16557, B1 => 
                           REGISTERS_10_3_port, B2 => n16560, ZN => n16492);
   U14714 : AOI22_X1 port map( A1 => REGISTERS_18_3_port, A2 => n16584, B1 => 
                           REGISTERS_21_3_port, B2 => n16568, ZN => n16491);
   U14715 : AOI22_X1 port map( A1 => REGISTERS_19_3_port, A2 => n16569, B1 => 
                           REGISTERS_17_3_port, B2 => n16579, ZN => n16490);
   U14716 : NAND4_X1 port map( A1 => n16493, A2 => n16492, A3 => n16491, A4 => 
                           n16490, ZN => n16494);
   U14717 : NOR3_X1 port map( A1 => n16496, A2 => n16495, A3 => n16494, ZN => 
                           n16502);
   U14718 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n16595, B1 => 
                           REGISTERS_7_3_port, B2 => n16454, ZN => n16500);
   U14719 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n16544, B1 => 
                           REGISTERS_5_3_port, B2 => n16518, ZN => n16499);
   U14720 : AOI22_X1 port map( A1 => REGISTERS_0_3_port, A2 => n16547, B1 => 
                           REGISTERS_2_3_port, B2 => n16596, ZN => n16498);
   U14721 : AOI22_X1 port map( A1 => REGISTERS_3_3_port, A2 => n16593, B1 => 
                           REGISTERS_6_3_port, B2 => n16546, ZN => n16497);
   U14722 : AND4_X1 port map( A1 => n16500, A2 => n16499, A3 => n16498, A4 => 
                           n16497, ZN => n16501);
   U14723 : OAI222_X1 port map( A1 => n15796, A2 => n16502, B1 => n16553, B2 =>
                           n16501, C1 => n16049, C2 => n8381, ZN => n8630);
   U14724 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n16562, B1 => 
                           REGISTERS_19_2_port, B2 => n16569, ZN => n16506);
   U14725 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n16557, B1 => 
                           REGISTERS_11_2_port, B2 => n15782, ZN => n16505);
   U14726 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n16559, B1 => 
                           REGISTERS_8_2_port, B2 => n16567, ZN => n16504);
   U14727 : AOI22_X1 port map( A1 => REGISTERS_18_2_port, A2 => n16584, B1 => 
                           REGISTERS_17_2_port, B2 => n16579, ZN => n16503);
   U14728 : NAND4_X1 port map( A1 => n16506, A2 => n16505, A3 => n16504, A4 => 
                           n16503, ZN => n16517);
   U14729 : AOI22_X1 port map( A1 => REGISTERS_15_2_port, A2 => n16558, B1 => 
                           REGISTERS_16_2_port, B2 => n16561, ZN => n16510);
   U14730 : AOI22_X1 port map( A1 => REGISTERS_31_2_port, A2 => n16583, B1 => 
                           REGISTERS_27_2_port, B2 => n16573, ZN => n16509);
   U14731 : AOI22_X1 port map( A1 => REGISTERS_14_2_port, A2 => n16571, B1 => 
                           REGISTERS_23_2_port, B2 => n16572, ZN => n16508);
   U14732 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n16570, B1 => 
                           REGISTERS_9_2_port, B2 => n16525, ZN => n16507);
   U14733 : NAND4_X1 port map( A1 => n16510, A2 => n16509, A3 => n16508, A4 => 
                           n16507, ZN => n16516);
   U14734 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n16581, B1 => 
                           REGISTERS_10_2_port, B2 => n16560, ZN => n16514);
   U14735 : AOI22_X1 port map( A1 => REGISTERS_26_2_port, A2 => n16582, B1 => 
                           REGISTERS_30_2_port, B2 => n16555, ZN => n16513);
   U14736 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n16568, B1 => 
                           REGISTERS_22_2_port, B2 => n16556, ZN => n16512);
   U14737 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n16580, B1 => 
                           REGISTERS_29_2_port, B2 => n16574, ZN => n16511);
   U14738 : NAND4_X1 port map( A1 => n16514, A2 => n16513, A3 => n16512, A4 => 
                           n16511, ZN => n16515);
   U14739 : NOR3_X1 port map( A1 => n16517, A2 => n16516, A3 => n16515, ZN => 
                           n16524);
   U14740 : AOI22_X1 port map( A1 => REGISTERS_0_2_port, A2 => n16597, B1 => 
                           REGISTERS_5_2_port, B2 => n16518, ZN => n16522);
   U14741 : AOI22_X1 port map( A1 => REGISTERS_6_2_port, A2 => n16592, B1 => 
                           REGISTERS_2_2_port, B2 => n16545, ZN => n16521);
   U14742 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n16595, B1 => 
                           REGISTERS_1_2_port, B2 => n16544, ZN => n16520);
   U14743 : AOI22_X1 port map( A1 => REGISTERS_3_2_port, A2 => n16593, B1 => 
                           REGISTERS_7_2_port, B2 => n16454, ZN => n16519);
   U14744 : AND4_X1 port map( A1 => n16522, A2 => n16521, A3 => n16520, A4 => 
                           n16519, ZN => n16523);
   U14745 : OAI222_X1 port map( A1 => n16605, A2 => n16524, B1 => n16603, B2 =>
                           n16523, C1 => n16071, C2 => n8380, ZN => n8631);
   U14746 : AOI22_X1 port map( A1 => REGISTERS_27_1_port, A2 => n16573, B1 => 
                           REGISTERS_12_1_port, B2 => n16580, ZN => n16529);
   U14747 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n16567, B1 => 
                           REGISTERS_22_1_port, B2 => n16556, ZN => n16528);
   U14748 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n16568, B1 => 
                           REGISTERS_17_1_port, B2 => n16579, ZN => n16527);
   U14749 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n16561, B1 => 
                           REGISTERS_9_1_port, B2 => n16525, ZN => n16526);
   U14750 : NAND4_X1 port map( A1 => n16529, A2 => n16528, A3 => n16527, A4 => 
                           n16526, ZN => n16541);
   U14751 : AOI22_X1 port map( A1 => REGISTERS_11_1_port, A2 => n16530, B1 => 
                           REGISTERS_10_1_port, B2 => n16560, ZN => n16534);
   U14752 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n16557, B1 => 
                           REGISTERS_30_1_port, B2 => n16555, ZN => n16533);
   U14753 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n16562, B1 => 
                           REGISTERS_15_1_port, B2 => n16558, ZN => n16532);
   U14754 : AOI22_X1 port map( A1 => REGISTERS_31_1_port, A2 => n16583, B1 => 
                           REGISTERS_26_1_port, B2 => n16582, ZN => n16531);
   U14755 : NAND4_X1 port map( A1 => n16534, A2 => n16533, A3 => n16532, A4 => 
                           n16531, ZN => n16540);
   U14756 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n16574, B1 => 
                           REGISTERS_23_1_port, B2 => n16572, ZN => n16538);
   U14757 : AOI22_X1 port map( A1 => REGISTERS_19_1_port, A2 => n16569, B1 => 
                           REGISTERS_28_1_port, B2 => n16570, ZN => n16537);
   U14758 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n16581, B1 => 
                           REGISTERS_14_1_port, B2 => n16571, ZN => n16536);
   U14759 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n16559, B1 => 
                           REGISTERS_18_1_port, B2 => n16584, ZN => n16535);
   U14760 : NAND4_X1 port map( A1 => n16538, A2 => n16537, A3 => n16536, A4 => 
                           n16535, ZN => n16539);
   U14761 : NOR3_X1 port map( A1 => n16541, A2 => n16540, A3 => n16539, ZN => 
                           n16554);
   U14762 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n16542, B1 => 
                           REGISTERS_7_1_port, B2 => n16454, ZN => n16551);
   U14763 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n16544, B1 => 
                           REGISTERS_4_1_port, B2 => n16543, ZN => n16550);
   U14764 : AOI22_X1 port map( A1 => REGISTERS_6_1_port, A2 => n16546, B1 => 
                           REGISTERS_2_1_port, B2 => n16545, ZN => n16549);
   U14765 : AOI22_X1 port map( A1 => REGISTERS_0_1_port, A2 => n16547, B1 => 
                           REGISTERS_3_1_port, B2 => n16593, ZN => n16548);
   U14766 : AND4_X1 port map( A1 => n16551, A2 => n16550, A3 => n16549, A4 => 
                           n16548, ZN => n16552);
   U14767 : OAI222_X1 port map( A1 => n15796, A2 => n16554, B1 => n16553, B2 =>
                           n16552, C1 => n16071, C2 => n8379, ZN => n8632);
   U14768 : AOI22_X1 port map( A1 => REGISTERS_22_0_port, A2 => n16556, B1 => 
                           REGISTERS_30_0_port, B2 => n16555, ZN => n16566);
   U14769 : AOI22_X1 port map( A1 => REGISTERS_15_0_port, A2 => n16558, B1 => 
                           REGISTERS_25_0_port, B2 => n16557, ZN => n16565);
   U14770 : AOI22_X1 port map( A1 => REGISTERS_10_0_port, A2 => n16560, B1 => 
                           REGISTERS_24_0_port, B2 => n16559, ZN => n16564);
   U14771 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n16562, B1 => 
                           REGISTERS_16_0_port, B2 => n16561, ZN => n16563);
   U14772 : NAND4_X1 port map( A1 => n16566, A2 => n16565, A3 => n16564, A4 => 
                           n16563, ZN => n16591);
   U14773 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n16568, B1 => 
                           REGISTERS_8_0_port, B2 => n16567, ZN => n16578);
   U14774 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n16570, B1 => 
                           REGISTERS_19_0_port, B2 => n16569, ZN => n16577);
   U14775 : AOI22_X1 port map( A1 => REGISTERS_23_0_port, A2 => n16572, B1 => 
                           REGISTERS_14_0_port, B2 => n16571, ZN => n16576);
   U14776 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n16574, B1 => 
                           REGISTERS_27_0_port, B2 => n16573, ZN => n16575);
   U14777 : NAND4_X1 port map( A1 => n16578, A2 => n16577, A3 => n16576, A4 => 
                           n16575, ZN => n16590);
   U14778 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n16579, B1 => 
                           REGISTERS_9_0_port, B2 => n16029, ZN => n16588);
   U14779 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n16581, B1 => 
                           REGISTERS_12_0_port, B2 => n16580, ZN => n16587);
   U14780 : AOI22_X1 port map( A1 => REGISTERS_31_0_port, A2 => n16583, B1 => 
                           REGISTERS_26_0_port, B2 => n16582, ZN => n16586);
   U14781 : AOI22_X1 port map( A1 => REGISTERS_18_0_port, A2 => n16584, B1 => 
                           REGISTERS_11_0_port, B2 => n16414, ZN => n16585);
   U14782 : NAND4_X1 port map( A1 => n16588, A2 => n16587, A3 => n16586, A4 => 
                           n16585, ZN => n16589);
   U14783 : NOR3_X1 port map( A1 => n16591, A2 => n16590, A3 => n16589, ZN => 
                           n16604);
   U14784 : AOI22_X1 port map( A1 => REGISTERS_6_0_port, A2 => n16592, B1 => 
                           REGISTERS_5_0_port, B2 => n16518, ZN => n16601);
   U14785 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n16544, B1 => 
                           REGISTERS_3_0_port, B2 => n16593, ZN => n16600);
   U14786 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n16595, B1 => 
                           REGISTERS_7_0_port, B2 => n16594, ZN => n16599);
   U14787 : AOI22_X1 port map( A1 => REGISTERS_0_0_port, A2 => n16597, B1 => 
                           REGISTERS_2_0_port, B2 => n16596, ZN => n16598);
   U14788 : OAI222_X1 port map( A1 => n16605, A2 => n16604, B1 => n16603, B2 =>
                           n16602, C1 => n16026, C2 => n8378, ZN => n8633);
   U14789 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1)
                           , ZN => n16714);
   U14790 : INV_X1 port map( A => ADD_WR(4), ZN => n16606);
   U14791 : NAND2_X1 port map( A1 => WR, A2 => n16606, ZN => n16644);
   U14792 : NAND2_X1 port map( A1 => n16714, A2 => n16639, ZN => n16610);
   U14793 : NAND2_X1 port map( A1 => n13731, A2 => n16608, ZN => n16609);
   U14794 : NAND2_X1 port map( A1 => DATAIN(63), A2 => n13731, ZN => n16745);
   U14795 : CLKBUF_X1 port map( A => n16745, Z => n16815);
   U14796 : OAI22_X1 port map( A1 => n16884, A2 => n16609, B1 => n16815, B2 => 
                           n16610, ZN => n4503);
   U14797 : CLKBUF_X2 port map( A => n16609, Z => n16607);
   U14798 : NAND2_X1 port map( A1 => DATAIN(62), A2 => n13731, ZN => n16746);
   U14799 : OAI22_X1 port map( A1 => n18017, A2 => n16607, B1 => n16608, B2 => 
                           n16746, ZN => n4502);
   U14800 : NAND2_X1 port map( A1 => DATAIN(61), A2 => n13731, ZN => n16747);
   U14801 : OAI22_X1 port map( A1 => n18243, A2 => n16609, B1 => n16610, B2 => 
                           n16747, ZN => n4501);
   U14802 : NAND2_X1 port map( A1 => DATAIN(60), A2 => n13731, ZN => n16748);
   U14803 : OAI22_X1 port map( A1 => n18018, A2 => n16607, B1 => n16610, B2 => 
                           n16748, ZN => n4500);
   U14804 : NAND2_X1 port map( A1 => DATAIN(59), A2 => n13731, ZN => n16749);
   U14805 : OAI22_X1 port map( A1 => n18244, A2 => n16607, B1 => n16610, B2 => 
                           n16749, ZN => n4499);
   U14806 : NAND2_X1 port map( A1 => DATAIN(58), A2 => n13731, ZN => n16750);
   U14807 : OAI22_X1 port map( A1 => n18019, A2 => n16607, B1 => n16610, B2 => 
                           n16750, ZN => n4498);
   U14808 : NAND2_X1 port map( A1 => DATAIN(57), A2 => n13731, ZN => n16751);
   U14809 : OAI22_X1 port map( A1 => n18020, A2 => n16607, B1 => n16608, B2 => 
                           n16751, ZN => n4497);
   U14810 : NAND2_X1 port map( A1 => DATAIN(56), A2 => n13731, ZN => n16752);
   U14811 : OAI22_X1 port map( A1 => n18245, A2 => n16607, B1 => n16610, B2 => 
                           n16752, ZN => n4496);
   U14812 : NAND2_X1 port map( A1 => DATAIN(55), A2 => n13731, ZN => n16753);
   U14813 : OAI22_X1 port map( A1 => n18246, A2 => n16607, B1 => n16610, B2 => 
                           n16753, ZN => n4495);
   U14814 : NAND2_X1 port map( A1 => DATAIN(54), A2 => n13731, ZN => n16754);
   U14815 : OAI22_X1 port map( A1 => n18021, A2 => n16607, B1 => n16610, B2 => 
                           n16754, ZN => n4494);
   U14816 : NAND2_X1 port map( A1 => DATAIN(53), A2 => n13731, ZN => n16755);
   U14817 : OAI22_X1 port map( A1 => n18247, A2 => n16607, B1 => n16608, B2 => 
                           n16755, ZN => n4493);
   U14818 : NAND2_X1 port map( A1 => DATAIN(52), A2 => n13731, ZN => n16756);
   U14819 : OAI22_X1 port map( A1 => n18248, A2 => n16607, B1 => n16610, B2 => 
                           n16756, ZN => n4492);
   U14820 : NAND2_X1 port map( A1 => DATAIN(51), A2 => n13731, ZN => n16757);
   U14821 : OAI22_X1 port map( A1 => n18022, A2 => n16609, B1 => n16608, B2 => 
                           n16757, ZN => n4491);
   U14822 : NAND2_X1 port map( A1 => DATAIN(50), A2 => n13731, ZN => n16758);
   U14823 : OAI22_X1 port map( A1 => n18023, A2 => n16607, B1 => n16608, B2 => 
                           n16758, ZN => n4490);
   U14824 : NAND2_X1 port map( A1 => DATAIN(49), A2 => n13731, ZN => n16759);
   U14825 : OAI22_X1 port map( A1 => n18024, A2 => n16607, B1 => n16610, B2 => 
                           n16759, ZN => n4489);
   U14826 : NAND2_X1 port map( A1 => DATAIN(48), A2 => n13731, ZN => n16760);
   U14827 : OAI22_X1 port map( A1 => n18249, A2 => n16609, B1 => n16610, B2 => 
                           n16760, ZN => n4488);
   U14828 : NAND2_X1 port map( A1 => DATAIN(47), A2 => n13731, ZN => n16761);
   U14829 : OAI22_X1 port map( A1 => n17388, A2 => n16609, B1 => n16608, B2 => 
                           n16761, ZN => n4487);
   U14830 : NAND2_X1 port map( A1 => DATAIN(46), A2 => n13731, ZN => n16762);
   U14831 : OAI22_X1 port map( A1 => n17172, A2 => n16607, B1 => n16608, B2 => 
                           n16762, ZN => n4486);
   U14832 : NAND2_X1 port map( A1 => DATAIN(45), A2 => n13731, ZN => n16763);
   U14833 : OAI22_X1 port map( A1 => n17389, A2 => n16607, B1 => n16608, B2 => 
                           n16763, ZN => n4485);
   U14834 : NAND2_X1 port map( A1 => DATAIN(44), A2 => n13731, ZN => n16764);
   U14835 : OAI22_X1 port map( A1 => n17173, A2 => n16609, B1 => n16608, B2 => 
                           n16764, ZN => n4484);
   U14836 : NAND2_X1 port map( A1 => DATAIN(43), A2 => n13731, ZN => n16765);
   U14837 : OAI22_X1 port map( A1 => n17390, A2 => n16609, B1 => n16608, B2 => 
                           n16765, ZN => n4483);
   U14838 : NAND2_X1 port map( A1 => DATAIN(42), A2 => n13731, ZN => n16766);
   U14839 : OAI22_X1 port map( A1 => n17174, A2 => n16607, B1 => n16608, B2 => 
                           n16766, ZN => n4482);
   U14840 : NAND2_X1 port map( A1 => DATAIN(41), A2 => n13731, ZN => n16767);
   U14841 : OAI22_X1 port map( A1 => n17175, A2 => n16607, B1 => n16608, B2 => 
                           n16767, ZN => n4481);
   U14842 : NAND2_X1 port map( A1 => DATAIN(40), A2 => n13731, ZN => n16768);
   U14843 : OAI22_X1 port map( A1 => n17176, A2 => n16607, B1 => n16608, B2 => 
                           n16768, ZN => n4480);
   U14844 : NAND2_X1 port map( A1 => DATAIN(39), A2 => n13731, ZN => n16769);
   U14845 : OAI22_X1 port map( A1 => n17177, A2 => n16607, B1 => n16608, B2 => 
                           n16769, ZN => n4479);
   U14846 : NAND2_X1 port map( A1 => DATAIN(38), A2 => n13731, ZN => n16770);
   U14847 : OAI22_X1 port map( A1 => n17178, A2 => n16609, B1 => n16608, B2 => 
                           n16770, ZN => n4478);
   U14848 : NAND2_X1 port map( A1 => DATAIN(37), A2 => n13731, ZN => n16771);
   U14849 : OAI22_X1 port map( A1 => n17179, A2 => n16607, B1 => n16608, B2 => 
                           n16771, ZN => n4477);
   U14850 : NAND2_X1 port map( A1 => DATAIN(36), A2 => n13731, ZN => n16772);
   U14851 : OAI22_X1 port map( A1 => n17391, A2 => n16609, B1 => n16608, B2 => 
                           n16772, ZN => n4476);
   U14852 : CLKBUF_X2 port map( A => n16610, Z => n16608);
   U14853 : NAND2_X1 port map( A1 => DATAIN(35), A2 => n13731, ZN => n16773);
   U14854 : OAI22_X1 port map( A1 => n18025, A2 => n16607, B1 => n16608, B2 => 
                           n16773, ZN => n4475);
   U14855 : NAND2_X1 port map( A1 => DATAIN(34), A2 => n13731, ZN => n16774);
   U14856 : OAI22_X1 port map( A1 => n18250, A2 => n16609, B1 => n16610, B2 => 
                           n16774, ZN => n4474);
   U14857 : NAND2_X1 port map( A1 => DATAIN(33), A2 => n13731, ZN => n16775);
   U14858 : OAI22_X1 port map( A1 => n18026, A2 => n16607, B1 => n16608, B2 => 
                           n16775, ZN => n4473);
   U14859 : NAND2_X1 port map( A1 => DATAIN(32), A2 => n13731, ZN => n16776);
   U14860 : OAI22_X1 port map( A1 => n18027, A2 => n16609, B1 => n16608, B2 => 
                           n16776, ZN => n4472);
   U14861 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n13731, ZN => n16777);
   U14862 : OAI22_X1 port map( A1 => n18251, A2 => n16607, B1 => n16610, B2 => 
                           n16777, ZN => n4471);
   U14863 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n13731, ZN => n16778);
   U14864 : OAI22_X1 port map( A1 => n18252, A2 => n16609, B1 => n16608, B2 => 
                           n16778, ZN => n4470);
   U14865 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n13731, ZN => n16779);
   U14866 : OAI22_X1 port map( A1 => n18253, A2 => n16607, B1 => n16610, B2 => 
                           n16779, ZN => n4469);
   U14867 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n13731, ZN => n16781);
   U14868 : OAI22_X1 port map( A1 => n18254, A2 => n16609, B1 => n16608, B2 => 
                           n16781, ZN => n4468);
   U14869 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n13731, ZN => n16782);
   U14870 : OAI22_X1 port map( A1 => n17180, A2 => n16609, B1 => n16610, B2 => 
                           n16782, ZN => n4467);
   U14871 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n13731, ZN => n16783);
   U14872 : OAI22_X1 port map( A1 => n17392, A2 => n16607, B1 => n16608, B2 => 
                           n16783, ZN => n4466);
   U14873 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n13731, ZN => n16784);
   U14874 : OAI22_X1 port map( A1 => n17393, A2 => n16609, B1 => n16610, B2 => 
                           n16784, ZN => n4465);
   U14875 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n13731, ZN => n16785);
   U14876 : OAI22_X1 port map( A1 => n17394, A2 => n16607, B1 => n16608, B2 => 
                           n16785, ZN => n4464);
   U14877 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n13731, ZN => n16786);
   U14878 : OAI22_X1 port map( A1 => n17181, A2 => n16609, B1 => n16610, B2 => 
                           n16786, ZN => n4463);
   U14879 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n13731, ZN => n16787);
   U14880 : OAI22_X1 port map( A1 => n17182, A2 => n16607, B1 => n16610, B2 => 
                           n16787, ZN => n4462);
   U14881 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n13731, ZN => n16788);
   U14882 : OAI22_X1 port map( A1 => n17395, A2 => n16607, B1 => n16608, B2 => 
                           n16788, ZN => n4461);
   U14883 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n13731, ZN => n16789);
   U14884 : OAI22_X1 port map( A1 => n17183, A2 => n16607, B1 => n16608, B2 => 
                           n16789, ZN => n4460);
   U14885 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n13731, ZN => n16790);
   U14886 : OAI22_X1 port map( A1 => n17184, A2 => n16607, B1 => n16610, B2 => 
                           n16790, ZN => n4459);
   U14887 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n13731, ZN => n16791);
   U14888 : OAI22_X1 port map( A1 => n17396, A2 => n16607, B1 => n16610, B2 => 
                           n16791, ZN => n4458);
   U14889 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n13731, ZN => n16792);
   U14890 : OAI22_X1 port map( A1 => n17185, A2 => n16607, B1 => n16608, B2 => 
                           n16792, ZN => n4457);
   U14891 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n13731, ZN => n16793);
   U14892 : OAI22_X1 port map( A1 => n17397, A2 => n16607, B1 => n16608, B2 => 
                           n16793, ZN => n4456);
   U14893 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n13731, ZN => n16794);
   U14894 : OAI22_X1 port map( A1 => n18028, A2 => n16609, B1 => n16610, B2 => 
                           n16794, ZN => n4455);
   U14895 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n13731, ZN => n16795);
   U14896 : OAI22_X1 port map( A1 => n18029, A2 => n16609, B1 => n16610, B2 => 
                           n16795, ZN => n4454);
   U14897 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n13731, ZN => n16796);
   U14898 : OAI22_X1 port map( A1 => n18255, A2 => n16607, B1 => n16608, B2 => 
                           n16796, ZN => n4453);
   U14899 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n13731, ZN => n16797);
   U14900 : OAI22_X1 port map( A1 => n17398, A2 => n16607, B1 => n16608, B2 => 
                           n16797, ZN => n4452);
   U14901 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n13731, ZN => n16798);
   U14902 : OAI22_X1 port map( A1 => n17399, A2 => n16609, B1 => n16608, B2 => 
                           n16798, ZN => n4451);
   U14903 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n13731, ZN => n16799);
   U14904 : OAI22_X1 port map( A1 => n17186, A2 => n16607, B1 => n16608, B2 => 
                           n16799, ZN => n4450);
   U14905 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n13731, ZN => n16800);
   U14906 : OAI22_X1 port map( A1 => n17187, A2 => n16609, B1 => n16608, B2 => 
                           n16800, ZN => n4449);
   U14907 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n13731, ZN => n16801);
   U14908 : OAI22_X1 port map( A1 => n17188, A2 => n16607, B1 => n16608, B2 => 
                           n16801, ZN => n4448);
   U14909 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n13731, ZN => n16802);
   U14910 : OAI22_X1 port map( A1 => n17400, A2 => n16609, B1 => n16608, B2 => 
                           n16802, ZN => n4447);
   U14911 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n13731, ZN => n16803);
   U14912 : OAI22_X1 port map( A1 => n17189, A2 => n16609, B1 => n16608, B2 => 
                           n16803, ZN => n4446);
   U14913 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n13731, ZN => n16804);
   U14914 : OAI22_X1 port map( A1 => n17401, A2 => n16607, B1 => n16608, B2 => 
                           n16804, ZN => n4445);
   U14915 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n13731, ZN => n16805);
   U14916 : OAI22_X1 port map( A1 => n17402, A2 => n16607, B1 => n16608, B2 => 
                           n16805, ZN => n4444);
   U14917 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n13731, ZN => n16806);
   U14918 : OAI22_X1 port map( A1 => n17403, A2 => n16609, B1 => n16608, B2 => 
                           n16806, ZN => n4443);
   U14919 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n13731, ZN => n16808);
   U14920 : OAI22_X1 port map( A1 => n17404, A2 => n16607, B1 => n16610, B2 => 
                           n16808, ZN => n4442);
   U14921 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n13731, ZN => n16810);
   U14922 : OAI22_X1 port map( A1 => n17405, A2 => n16609, B1 => n16608, B2 => 
                           n16810, ZN => n4441);
   U14923 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n13731, ZN => n16812);
   U14924 : OAI22_X1 port map( A1 => n18256, A2 => n16607, B1 => n16610, B2 => 
                           n16812, ZN => n4440);
   U14925 : INV_X1 port map( A => ADD_WR(0), ZN => n16627);
   U14926 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n16627, 
                           ZN => n16719);
   U14927 : NAND2_X1 port map( A1 => n16639, A2 => n16719, ZN => n16612);
   U14928 : CLKBUF_X2 port map( A => n16612, Z => n16614);
   U14929 : NAND2_X1 port map( A1 => n13731, A2 => n16614, ZN => n16613);
   U14930 : OAI22_X1 port map( A1 => n17105, A2 => n16613, B1 => n16745, B2 => 
                           n16614, ZN => n4439);
   U14931 : CLKBUF_X2 port map( A => n16613, Z => n16611);
   U14932 : CLKBUF_X1 port map( A => n16746, Z => n16816);
   U14933 : OAI22_X1 port map( A1 => n18257, A2 => n16611, B1 => n16816, B2 => 
                           n16612, ZN => n4438);
   U14934 : CLKBUF_X1 port map( A => n16747, Z => n16817);
   U14935 : OAI22_X1 port map( A1 => n18701, A2 => n16613, B1 => n16817, B2 => 
                           n16614, ZN => n4437);
   U14936 : CLKBUF_X1 port map( A => n16748, Z => n16818);
   U14937 : OAI22_X1 port map( A1 => n18258, A2 => n16611, B1 => n16818, B2 => 
                           n16612, ZN => n4436);
   U14938 : CLKBUF_X1 port map( A => n16749, Z => n16819);
   U14939 : OAI22_X1 port map( A1 => n18702, A2 => n16611, B1 => n16819, B2 => 
                           n16612, ZN => n4435);
   U14940 : CLKBUF_X1 port map( A => n16750, Z => n16820);
   U14941 : OAI22_X1 port map( A1 => n18259, A2 => n16611, B1 => n16820, B2 => 
                           n16614, ZN => n4434);
   U14942 : CLKBUF_X1 port map( A => n16751, Z => n16821);
   U14943 : OAI22_X1 port map( A1 => n18703, A2 => n16611, B1 => n16821, B2 => 
                           n16612, ZN => n4433);
   U14944 : OAI22_X1 port map( A1 => n18260, A2 => n16611, B1 => n16822, B2 => 
                           n16614, ZN => n4432);
   U14945 : CLKBUF_X1 port map( A => n16753, Z => n16823);
   U14946 : OAI22_X1 port map( A1 => n18030, A2 => n16611, B1 => n16823, B2 => 
                           n16614, ZN => n4431);
   U14947 : CLKBUF_X1 port map( A => n16754, Z => n16824);
   U14948 : OAI22_X1 port map( A1 => n18704, A2 => n16611, B1 => n16824, B2 => 
                           n16614, ZN => n4430);
   U14949 : CLKBUF_X1 port map( A => n16755, Z => n16825);
   U14950 : OAI22_X1 port map( A1 => n18261, A2 => n16611, B1 => n16825, B2 => 
                           n16614, ZN => n4429);
   U14951 : CLKBUF_X1 port map( A => n16756, Z => n16826);
   U14952 : OAI22_X1 port map( A1 => n18262, A2 => n16611, B1 => n16826, B2 => 
                           n16614, ZN => n4428);
   U14953 : CLKBUF_X1 port map( A => n16757, Z => n16827);
   U14954 : OAI22_X1 port map( A1 => n18263, A2 => n16613, B1 => n16827, B2 => 
                           n16612, ZN => n4427);
   U14955 : CLKBUF_X1 port map( A => n16758, Z => n16828);
   U14956 : OAI22_X1 port map( A1 => n18705, A2 => n16611, B1 => n16828, B2 => 
                           n16612, ZN => n4426);
   U14957 : CLKBUF_X1 port map( A => n16759, Z => n16829);
   U14958 : OAI22_X1 port map( A1 => n18706, A2 => n16611, B1 => n16829, B2 => 
                           n16612, ZN => n4425);
   U14959 : CLKBUF_X1 port map( A => n16760, Z => n16830);
   U14960 : OAI22_X1 port map( A1 => n18707, A2 => n16613, B1 => n16830, B2 => 
                           n16614, ZN => n4424);
   U14961 : CLKBUF_X1 port map( A => n16761, Z => n16831);
   U14962 : OAI22_X1 port map( A1 => n18264, A2 => n16613, B1 => n16831, B2 => 
                           n16612, ZN => n4423);
   U14963 : CLKBUF_X1 port map( A => n16762, Z => n16832);
   U14964 : OAI22_X1 port map( A1 => n18265, A2 => n16611, B1 => n16832, B2 => 
                           n16612, ZN => n4422);
   U14965 : CLKBUF_X1 port map( A => n16763, Z => n16833);
   U14966 : OAI22_X1 port map( A1 => n18708, A2 => n16611, B1 => n16833, B2 => 
                           n16612, ZN => n4421);
   U14967 : CLKBUF_X1 port map( A => n16764, Z => n16834);
   U14968 : OAI22_X1 port map( A1 => n18266, A2 => n16613, B1 => n16834, B2 => 
                           n16614, ZN => n4420);
   U14969 : CLKBUF_X1 port map( A => n16765, Z => n16835);
   U14970 : OAI22_X1 port map( A1 => n18267, A2 => n16613, B1 => n16835, B2 => 
                           n16612, ZN => n4419);
   U14971 : CLKBUF_X1 port map( A => n16766, Z => n16836);
   U14972 : OAI22_X1 port map( A1 => n18709, A2 => n16611, B1 => n16836, B2 => 
                           n16614, ZN => n4418);
   U14973 : OAI22_X1 port map( A1 => n18268, A2 => n16611, B1 => n16837, B2 => 
                           n16614, ZN => n4417);
   U14974 : CLKBUF_X1 port map( A => n16768, Z => n16838);
   U14975 : OAI22_X1 port map( A1 => n18031, A2 => n16611, B1 => n16838, B2 => 
                           n16612, ZN => n4416);
   U14976 : CLKBUF_X1 port map( A => n16769, Z => n16839);
   U14977 : OAI22_X1 port map( A1 => n18269, A2 => n16611, B1 => n16839, B2 => 
                           n16614, ZN => n4415);
   U14978 : CLKBUF_X1 port map( A => n16770, Z => n16840);
   U14979 : OAI22_X1 port map( A1 => n18270, A2 => n16613, B1 => n16840, B2 => 
                           n16612, ZN => n4414);
   U14980 : CLKBUF_X1 port map( A => n16771, Z => n16841);
   U14981 : OAI22_X1 port map( A1 => n18271, A2 => n16611, B1 => n16841, B2 => 
                           n16612, ZN => n4413);
   U14982 : CLKBUF_X1 port map( A => n16772, Z => n16842);
   U14983 : OAI22_X1 port map( A1 => n18272, A2 => n16613, B1 => n16842, B2 => 
                           n16612, ZN => n4412);
   U14984 : CLKBUF_X1 port map( A => n16773, Z => n16843);
   U14985 : OAI22_X1 port map( A1 => n18710, A2 => n16611, B1 => n16843, B2 => 
                           n16612, ZN => n4411);
   U14986 : CLKBUF_X1 port map( A => n16774, Z => n16844);
   U14987 : OAI22_X1 port map( A1 => n18273, A2 => n16613, B1 => n16844, B2 => 
                           n16612, ZN => n4410);
   U14988 : CLKBUF_X1 port map( A => n16775, Z => n16845);
   U14989 : OAI22_X1 port map( A1 => n18274, A2 => n16611, B1 => n16845, B2 => 
                           n16612, ZN => n4409);
   U14990 : CLKBUF_X1 port map( A => n16776, Z => n16846);
   U14991 : OAI22_X1 port map( A1 => n18275, A2 => n16613, B1 => n16846, B2 => 
                           n16612, ZN => n4408);
   U14992 : CLKBUF_X1 port map( A => n16777, Z => n16847);
   U14993 : OAI22_X1 port map( A1 => n18032, A2 => n16611, B1 => n16847, B2 => 
                           n16612, ZN => n4407);
   U14994 : CLKBUF_X1 port map( A => n16778, Z => n16848);
   U14995 : OAI22_X1 port map( A1 => n18711, A2 => n16613, B1 => n16848, B2 => 
                           n16612, ZN => n4406);
   U14996 : CLKBUF_X1 port map( A => n16779, Z => n16849);
   U14997 : OAI22_X1 port map( A1 => n18276, A2 => n16611, B1 => n16849, B2 => 
                           n16612, ZN => n4405);
   U14998 : CLKBUF_X1 port map( A => n16781, Z => n16850);
   U14999 : OAI22_X1 port map( A1 => n18277, A2 => n16613, B1 => n16850, B2 => 
                           n16614, ZN => n4404);
   U15000 : OAI22_X1 port map( A1 => n17794, A2 => n16613, B1 => n16851, B2 => 
                           n16614, ZN => n4403);
   U15001 : CLKBUF_X1 port map( A => n16783, Z => n16852);
   U15002 : OAI22_X1 port map( A1 => n17406, A2 => n16611, B1 => n16852, B2 => 
                           n16614, ZN => n4402);
   U15003 : CLKBUF_X1 port map( A => n16784, Z => n16853);
   U15004 : OAI22_X1 port map( A1 => n17795, A2 => n16613, B1 => n16853, B2 => 
                           n16614, ZN => n4401);
   U15005 : CLKBUF_X1 port map( A => n16785, Z => n16854);
   U15006 : OAI22_X1 port map( A1 => n17407, A2 => n16611, B1 => n16854, B2 => 
                           n16614, ZN => n4400);
   U15007 : CLKBUF_X1 port map( A => n16786, Z => n16855);
   U15008 : OAI22_X1 port map( A1 => n17796, A2 => n16613, B1 => n16855, B2 => 
                           n16614, ZN => n4399);
   U15009 : CLKBUF_X1 port map( A => n16787, Z => n16856);
   U15010 : OAI22_X1 port map( A1 => n17408, A2 => n16611, B1 => n16856, B2 => 
                           n16614, ZN => n4398);
   U15011 : CLKBUF_X1 port map( A => n16788, Z => n16857);
   U15012 : OAI22_X1 port map( A1 => n17190, A2 => n16611, B1 => n16857, B2 => 
                           n16614, ZN => n4397);
   U15013 : CLKBUF_X1 port map( A => n16789, Z => n16858);
   U15014 : OAI22_X1 port map( A1 => n17191, A2 => n16611, B1 => n16858, B2 => 
                           n16614, ZN => n4396);
   U15015 : CLKBUF_X1 port map( A => n16790, Z => n16859);
   U15016 : OAI22_X1 port map( A1 => n17409, A2 => n16611, B1 => n16859, B2 => 
                           n16614, ZN => n4395);
   U15017 : CLKBUF_X1 port map( A => n16791, Z => n16860);
   U15018 : OAI22_X1 port map( A1 => n17797, A2 => n16611, B1 => n16860, B2 => 
                           n16614, ZN => n4394);
   U15019 : CLKBUF_X1 port map( A => n16792, Z => n16861);
   U15020 : OAI22_X1 port map( A1 => n17798, A2 => n16611, B1 => n16861, B2 => 
                           n16614, ZN => n4393);
   U15021 : CLKBUF_X1 port map( A => n16793, Z => n16862);
   U15022 : OAI22_X1 port map( A1 => n17799, A2 => n16611, B1 => n16862, B2 => 
                           n16614, ZN => n4392);
   U15023 : CLKBUF_X1 port map( A => n16794, Z => n16863);
   U15024 : OAI22_X1 port map( A1 => n18712, A2 => n16613, B1 => n16863, B2 => 
                           n16614, ZN => n4391);
   U15025 : CLKBUF_X1 port map( A => n16795, Z => n16864);
   U15026 : OAI22_X1 port map( A1 => n18713, A2 => n16613, B1 => n16864, B2 => 
                           n16614, ZN => n4390);
   U15027 : CLKBUF_X1 port map( A => n16796, Z => n16865);
   U15028 : OAI22_X1 port map( A1 => n18714, A2 => n16611, B1 => n16865, B2 => 
                           n16614, ZN => n4389);
   U15029 : OAI22_X1 port map( A1 => n18278, A2 => n16611, B1 => n16866, B2 => 
                           n16614, ZN => n4388);
   U15030 : CLKBUF_X1 port map( A => n16798, Z => n16867);
   U15031 : OAI22_X1 port map( A1 => n18715, A2 => n16613, B1 => n16867, B2 => 
                           n16614, ZN => n4387);
   U15032 : CLKBUF_X1 port map( A => n16799, Z => n16868);
   U15033 : OAI22_X1 port map( A1 => n18033, A2 => n16611, B1 => n16868, B2 => 
                           n16614, ZN => n4386);
   U15034 : CLKBUF_X1 port map( A => n16800, Z => n16869);
   U15035 : OAI22_X1 port map( A1 => n18279, A2 => n16613, B1 => n16869, B2 => 
                           n16614, ZN => n4385);
   U15036 : CLKBUF_X1 port map( A => n16801, Z => n16870);
   U15037 : OAI22_X1 port map( A1 => n18280, A2 => n16611, B1 => n16870, B2 => 
                           n16614, ZN => n4384);
   U15038 : CLKBUF_X1 port map( A => n16802, Z => n16871);
   U15039 : OAI22_X1 port map( A1 => n18281, A2 => n16613, B1 => n16871, B2 => 
                           n16614, ZN => n4383);
   U15040 : CLKBUF_X1 port map( A => n16803, Z => n16872);
   U15041 : OAI22_X1 port map( A1 => n18282, A2 => n16613, B1 => n16872, B2 => 
                           n16614, ZN => n4382);
   U15042 : CLKBUF_X1 port map( A => n16804, Z => n16873);
   U15043 : OAI22_X1 port map( A1 => n18283, A2 => n16611, B1 => n16873, B2 => 
                           n16614, ZN => n4381);
   U15044 : CLKBUF_X1 port map( A => n16805, Z => n16874);
   U15045 : OAI22_X1 port map( A1 => n18716, A2 => n16611, B1 => n16874, B2 => 
                           n16612, ZN => n4380);
   U15046 : CLKBUF_X1 port map( A => n16806, Z => n16875);
   U15047 : OAI22_X1 port map( A1 => n18717, A2 => n16613, B1 => n16875, B2 => 
                           n16614, ZN => n4379);
   U15048 : CLKBUF_X1 port map( A => n16808, Z => n16876);
   U15049 : OAI22_X1 port map( A1 => n18284, A2 => n16611, B1 => n16876, B2 => 
                           n16614, ZN => n4378);
   U15050 : CLKBUF_X1 port map( A => n16810, Z => n16878);
   U15051 : OAI22_X1 port map( A1 => n18718, A2 => n16613, B1 => n16878, B2 => 
                           n16612, ZN => n4377);
   U15052 : CLKBUF_X1 port map( A => n16812, Z => n16881);
   U15053 : OAI22_X1 port map( A1 => n18719, A2 => n16611, B1 => n16881, B2 => 
                           n16614, ZN => n4376);
   U15054 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n16627, ZN => n16632);
   U15055 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n16632, ZN => n16724);
   U15056 : NAND2_X1 port map( A1 => n16639, A2 => n16724, ZN => n16615);
   U15057 : CLKBUF_X2 port map( A => n16615, Z => n16617);
   U15058 : NAND2_X1 port map( A1 => n13731, A2 => n16617, ZN => n16616);
   U15059 : OAI22_X1 port map( A1 => n17106, A2 => n16616, B1 => n16815, B2 => 
                           n16617, ZN => n4375);
   U15060 : OAI22_X1 port map( A1 => n18720, A2 => n16618, B1 => n16746, B2 => 
                           n16615, ZN => n4374);
   U15061 : OAI22_X1 port map( A1 => n18285, A2 => n16616, B1 => n16747, B2 => 
                           n16617, ZN => n4373);
   U15062 : OAI22_X1 port map( A1 => n18721, A2 => n16618, B1 => n16748, B2 => 
                           n16615, ZN => n4372);
   U15063 : OAI22_X1 port map( A1 => n18722, A2 => n16618, B1 => n16749, B2 => 
                           n16615, ZN => n4371);
   U15064 : OAI22_X1 port map( A1 => n18723, A2 => n16616, B1 => n16750, B2 => 
                           n16617, ZN => n4370);
   U15065 : OAI22_X1 port map( A1 => n18286, A2 => n16618, B1 => n16751, B2 => 
                           n16615, ZN => n4369);
   U15066 : OAI22_X1 port map( A1 => n18287, A2 => n16616, B1 => n16752, B2 => 
                           n16617, ZN => n4368);
   U15067 : OAI22_X1 port map( A1 => n18288, A2 => n16618, B1 => n16753, B2 => 
                           n16617, ZN => n4367);
   U15068 : OAI22_X1 port map( A1 => n18724, A2 => n16616, B1 => n16754, B2 => 
                           n16617, ZN => n4366);
   U15069 : OAI22_X1 port map( A1 => n18725, A2 => n16618, B1 => n16755, B2 => 
                           n16617, ZN => n4365);
   U15070 : OAI22_X1 port map( A1 => n18289, A2 => n16618, B1 => n16756, B2 => 
                           n16617, ZN => n4364);
   U15071 : OAI22_X1 port map( A1 => n18726, A2 => n16616, B1 => n16757, B2 => 
                           n16615, ZN => n4363);
   U15072 : OAI22_X1 port map( A1 => n18727, A2 => n16618, B1 => n16758, B2 => 
                           n16615, ZN => n4362);
   U15073 : OAI22_X1 port map( A1 => n18290, A2 => n16618, B1 => n16759, B2 => 
                           n16615, ZN => n4361);
   U15074 : OAI22_X1 port map( A1 => n18728, A2 => n16616, B1 => n16760, B2 => 
                           n16617, ZN => n4360);
   U15075 : OAI22_X1 port map( A1 => n18291, A2 => n16616, B1 => n16761, B2 => 
                           n16615, ZN => n4359);
   U15076 : OAI22_X1 port map( A1 => n18729, A2 => n16618, B1 => n16762, B2 => 
                           n16615, ZN => n4358);
   U15077 : OAI22_X1 port map( A1 => n18730, A2 => n16618, B1 => n16763, B2 => 
                           n16615, ZN => n4357);
   U15078 : OAI22_X1 port map( A1 => n18731, A2 => n16616, B1 => n16764, B2 => 
                           n16617, ZN => n4356);
   U15079 : OAI22_X1 port map( A1 => n18732, A2 => n16616, B1 => n16765, B2 => 
                           n16615, ZN => n4355);
   U15080 : OAI22_X1 port map( A1 => n18292, A2 => n16618, B1 => n16766, B2 => 
                           n16617, ZN => n4354);
   U15081 : OAI22_X1 port map( A1 => n18293, A2 => n16618, B1 => n16767, B2 => 
                           n16617, ZN => n4353);
   U15082 : OAI22_X1 port map( A1 => n18733, A2 => n16618, B1 => n16768, B2 => 
                           n16615, ZN => n4352);
   U15083 : OAI22_X1 port map( A1 => n18734, A2 => n16618, B1 => n16769, B2 => 
                           n16617, ZN => n4351);
   U15084 : OAI22_X1 port map( A1 => n18735, A2 => n16616, B1 => n16770, B2 => 
                           n16615, ZN => n4350);
   U15085 : OAI22_X1 port map( A1 => n18736, A2 => n16618, B1 => n16771, B2 => 
                           n16615, ZN => n4349);
   U15086 : OAI22_X1 port map( A1 => n18294, A2 => n16616, B1 => n16772, B2 => 
                           n16615, ZN => n4348);
   U15087 : OAI22_X1 port map( A1 => n18295, A2 => n16618, B1 => n16773, B2 => 
                           n16615, ZN => n4347);
   U15088 : OAI22_X1 port map( A1 => n18737, A2 => n16616, B1 => n16774, B2 => 
                           n16615, ZN => n4346);
   U15089 : OAI22_X1 port map( A1 => n18738, A2 => n16618, B1 => n16775, B2 => 
                           n16615, ZN => n4345);
   U15090 : OAI22_X1 port map( A1 => n18296, A2 => n16616, B1 => n16776, B2 => 
                           n16615, ZN => n4344);
   U15091 : OAI22_X1 port map( A1 => n18297, A2 => n16618, B1 => n16777, B2 => 
                           n16615, ZN => n4343);
   U15092 : OAI22_X1 port map( A1 => n18298, A2 => n16616, B1 => n16778, B2 => 
                           n16615, ZN => n4342);
   U15093 : OAI22_X1 port map( A1 => n18299, A2 => n16618, B1 => n16779, B2 => 
                           n16615, ZN => n4341);
   U15094 : OAI22_X1 port map( A1 => n18300, A2 => n16616, B1 => n16781, B2 => 
                           n16617, ZN => n4340);
   U15095 : CLKBUF_X2 port map( A => n16616, Z => n16618);
   U15096 : OAI22_X1 port map( A1 => n17800, A2 => n16618, B1 => n16782, B2 => 
                           n16617, ZN => n4339);
   U15097 : OAI22_X1 port map( A1 => n17801, A2 => n16618, B1 => n16783, B2 => 
                           n16617, ZN => n4338);
   U15098 : OAI22_X1 port map( A1 => n17410, A2 => n16618, B1 => n16784, B2 => 
                           n16617, ZN => n4337);
   U15099 : OAI22_X1 port map( A1 => n17411, A2 => n16618, B1 => n16785, B2 => 
                           n16617, ZN => n4336);
   U15100 : OAI22_X1 port map( A1 => n17412, A2 => n16618, B1 => n16786, B2 => 
                           n16617, ZN => n4335);
   U15101 : OAI22_X1 port map( A1 => n17802, A2 => n16618, B1 => n16787, B2 => 
                           n16617, ZN => n4334);
   U15102 : OAI22_X1 port map( A1 => n17803, A2 => n16618, B1 => n16788, B2 => 
                           n16617, ZN => n4333);
   U15103 : OAI22_X1 port map( A1 => n17804, A2 => n16618, B1 => n16789, B2 => 
                           n16617, ZN => n4332);
   U15104 : OAI22_X1 port map( A1 => n17805, A2 => n16618, B1 => n16790, B2 => 
                           n16617, ZN => n4331);
   U15105 : OAI22_X1 port map( A1 => n17806, A2 => n16618, B1 => n16791, B2 => 
                           n16617, ZN => n4330);
   U15106 : OAI22_X1 port map( A1 => n17413, A2 => n16618, B1 => n16792, B2 => 
                           n16617, ZN => n4329);
   U15107 : OAI22_X1 port map( A1 => n17414, A2 => n16618, B1 => n16793, B2 => 
                           n16617, ZN => n4328);
   U15108 : OAI22_X1 port map( A1 => n18301, A2 => n16616, B1 => n16794, B2 => 
                           n16617, ZN => n4327);
   U15109 : OAI22_X1 port map( A1 => n18739, A2 => n16616, B1 => n16795, B2 => 
                           n16617, ZN => n4326);
   U15110 : OAI22_X1 port map( A1 => n18302, A2 => n16618, B1 => n16796, B2 => 
                           n16617, ZN => n4325);
   U15111 : OAI22_X1 port map( A1 => n18303, A2 => n16618, B1 => n16797, B2 => 
                           n16617, ZN => n4324);
   U15112 : OAI22_X1 port map( A1 => n18740, A2 => n16616, B1 => n16798, B2 => 
                           n16617, ZN => n4323);
   U15113 : OAI22_X1 port map( A1 => n18304, A2 => n16618, B1 => n16799, B2 => 
                           n16617, ZN => n4322);
   U15114 : OAI22_X1 port map( A1 => n18741, A2 => n16616, B1 => n16800, B2 => 
                           n16617, ZN => n4321);
   U15115 : OAI22_X1 port map( A1 => n18742, A2 => n16618, B1 => n16801, B2 => 
                           n16617, ZN => n4320);
   U15116 : OAI22_X1 port map( A1 => n18305, A2 => n16616, B1 => n16802, B2 => 
                           n16617, ZN => n4319);
   U15117 : OAI22_X1 port map( A1 => n18743, A2 => n16616, B1 => n16803, B2 => 
                           n16617, ZN => n4318);
   U15118 : OAI22_X1 port map( A1 => n18306, A2 => n16618, B1 => n16804, B2 => 
                           n16617, ZN => n4317);
   U15119 : OAI22_X1 port map( A1 => n18744, A2 => n16618, B1 => n16805, B2 => 
                           n16615, ZN => n4316);
   U15120 : OAI22_X1 port map( A1 => n18307, A2 => n16616, B1 => n16806, B2 => 
                           n16617, ZN => n4315);
   U15121 : OAI22_X1 port map( A1 => n18308, A2 => n16618, B1 => n16808, B2 => 
                           n16617, ZN => n4314);
   U15122 : OAI22_X1 port map( A1 => n18309, A2 => n16616, B1 => n16810, B2 => 
                           n16615, ZN => n4313);
   U15123 : OAI22_X1 port map( A1 => n18310, A2 => n16618, B1 => n16812, B2 => 
                           n16617, ZN => n4312);
   U15124 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n16637);
   U15125 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n16637, ZN => n16729);
   U15126 : NAND2_X1 port map( A1 => n16639, A2 => n16729, ZN => n16620);
   U15127 : CLKBUF_X2 port map( A => n16620, Z => n16622);
   U15128 : NAND2_X1 port map( A1 => n13731, A2 => n16622, ZN => n16621);
   U15129 : OAI22_X1 port map( A1 => n16963, A2 => n16621, B1 => n16745, B2 => 
                           n16622, ZN => n4311);
   U15130 : CLKBUF_X2 port map( A => n16621, Z => n16619);
   U15131 : OAI22_X1 port map( A1 => n18311, A2 => n16619, B1 => n16816, B2 => 
                           n16620, ZN => n4310);
   U15132 : OAI22_X1 port map( A1 => n18034, A2 => n16621, B1 => n16817, B2 => 
                           n16622, ZN => n4309);
   U15133 : OAI22_X1 port map( A1 => n18312, A2 => n16619, B1 => n16818, B2 => 
                           n16620, ZN => n4308);
   U15134 : OAI22_X1 port map( A1 => n18313, A2 => n16619, B1 => n16819, B2 => 
                           n16620, ZN => n4307);
   U15135 : OAI22_X1 port map( A1 => n18314, A2 => n16619, B1 => n16820, B2 => 
                           n16622, ZN => n4306);
   U15136 : OAI22_X1 port map( A1 => n18315, A2 => n16619, B1 => n16821, B2 => 
                           n16620, ZN => n4305);
   U15137 : OAI22_X1 port map( A1 => n18035, A2 => n16619, B1 => n16822, B2 => 
                           n16622, ZN => n4304);
   U15138 : OAI22_X1 port map( A1 => n18745, A2 => n16619, B1 => n16823, B2 => 
                           n16622, ZN => n4303);
   U15139 : OAI22_X1 port map( A1 => n18316, A2 => n16619, B1 => n16824, B2 => 
                           n16622, ZN => n4302);
   U15140 : OAI22_X1 port map( A1 => n18317, A2 => n16619, B1 => n16825, B2 => 
                           n16622, ZN => n4301);
   U15141 : OAI22_X1 port map( A1 => n18746, A2 => n16619, B1 => n16826, B2 => 
                           n16622, ZN => n4300);
   U15142 : OAI22_X1 port map( A1 => n18747, A2 => n16621, B1 => n16827, B2 => 
                           n16620, ZN => n4299);
   U15143 : OAI22_X1 port map( A1 => n18318, A2 => n16619, B1 => n16828, B2 => 
                           n16620, ZN => n4298);
   U15144 : OAI22_X1 port map( A1 => n18319, A2 => n16619, B1 => n16829, B2 => 
                           n16620, ZN => n4297);
   U15145 : OAI22_X1 port map( A1 => n18036, A2 => n16621, B1 => n16830, B2 => 
                           n16622, ZN => n4296);
   U15146 : OAI22_X1 port map( A1 => n18320, A2 => n16621, B1 => n16831, B2 => 
                           n16620, ZN => n4295);
   U15147 : OAI22_X1 port map( A1 => n18321, A2 => n16619, B1 => n16832, B2 => 
                           n16620, ZN => n4294);
   U15148 : OAI22_X1 port map( A1 => n18322, A2 => n16619, B1 => n16833, B2 => 
                           n16620, ZN => n4293);
   U15149 : OAI22_X1 port map( A1 => n18323, A2 => n16621, B1 => n16834, B2 => 
                           n16622, ZN => n4292);
   U15150 : OAI22_X1 port map( A1 => n18324, A2 => n16621, B1 => n16835, B2 => 
                           n16620, ZN => n4291);
   U15151 : OAI22_X1 port map( A1 => n18325, A2 => n16619, B1 => n16836, B2 => 
                           n16622, ZN => n4290);
   U15152 : OAI22_X1 port map( A1 => n18326, A2 => n16619, B1 => n16837, B2 => 
                           n16622, ZN => n4289);
   U15153 : OAI22_X1 port map( A1 => n18327, A2 => n16619, B1 => n16838, B2 => 
                           n16620, ZN => n4288);
   U15154 : OAI22_X1 port map( A1 => n18328, A2 => n16619, B1 => n16839, B2 => 
                           n16622, ZN => n4287);
   U15155 : OAI22_X1 port map( A1 => n18748, A2 => n16621, B1 => n16840, B2 => 
                           n16620, ZN => n4286);
   U15156 : OAI22_X1 port map( A1 => n18329, A2 => n16619, B1 => n16841, B2 => 
                           n16620, ZN => n4285);
   U15157 : OAI22_X1 port map( A1 => n18749, A2 => n16621, B1 => n16842, B2 => 
                           n16620, ZN => n4284);
   U15158 : OAI22_X1 port map( A1 => n18750, A2 => n16619, B1 => n16843, B2 => 
                           n16620, ZN => n4283);
   U15159 : OAI22_X1 port map( A1 => n18330, A2 => n16621, B1 => n16844, B2 => 
                           n16620, ZN => n4282);
   U15160 : OAI22_X1 port map( A1 => n18037, A2 => n16619, B1 => n16845, B2 => 
                           n16620, ZN => n4281);
   U15161 : OAI22_X1 port map( A1 => n18751, A2 => n16621, B1 => n16846, B2 => 
                           n16620, ZN => n4280);
   U15162 : OAI22_X1 port map( A1 => n18331, A2 => n16619, B1 => n16847, B2 => 
                           n16620, ZN => n4279);
   U15163 : OAI22_X1 port map( A1 => n18332, A2 => n16621, B1 => n16848, B2 => 
                           n16620, ZN => n4278);
   U15164 : OAI22_X1 port map( A1 => n18752, A2 => n16619, B1 => n16849, B2 => 
                           n16620, ZN => n4277);
   U15165 : OAI22_X1 port map( A1 => n18753, A2 => n16621, B1 => n16850, B2 => 
                           n16622, ZN => n4276);
   U15166 : OAI22_X1 port map( A1 => n17415, A2 => n16621, B1 => n16851, B2 => 
                           n16622, ZN => n4275);
   U15167 : OAI22_X1 port map( A1 => n17416, A2 => n16619, B1 => n16852, B2 => 
                           n16622, ZN => n4274);
   U15168 : OAI22_X1 port map( A1 => n17192, A2 => n16621, B1 => n16853, B2 => 
                           n16622, ZN => n4273);
   U15169 : OAI22_X1 port map( A1 => n17807, A2 => n16619, B1 => n16854, B2 => 
                           n16622, ZN => n4272);
   U15170 : OAI22_X1 port map( A1 => n17808, A2 => n16621, B1 => n16855, B2 => 
                           n16622, ZN => n4271);
   U15171 : OAI22_X1 port map( A1 => n17417, A2 => n16619, B1 => n16856, B2 => 
                           n16622, ZN => n4270);
   U15172 : OAI22_X1 port map( A1 => n17418, A2 => n16619, B1 => n16857, B2 => 
                           n16622, ZN => n4269);
   U15173 : OAI22_X1 port map( A1 => n17193, A2 => n16619, B1 => n16858, B2 => 
                           n16622, ZN => n4268);
   U15174 : OAI22_X1 port map( A1 => n17419, A2 => n16619, B1 => n16859, B2 => 
                           n16622, ZN => n4267);
   U15175 : OAI22_X1 port map( A1 => n17420, A2 => n16619, B1 => n16860, B2 => 
                           n16622, ZN => n4266);
   U15176 : OAI22_X1 port map( A1 => n17809, A2 => n16619, B1 => n16861, B2 => 
                           n16622, ZN => n4265);
   U15177 : OAI22_X1 port map( A1 => n17421, A2 => n16619, B1 => n16862, B2 => 
                           n16622, ZN => n4264);
   U15178 : OAI22_X1 port map( A1 => n18754, A2 => n16621, B1 => n16863, B2 => 
                           n16622, ZN => n4263);
   U15179 : OAI22_X1 port map( A1 => n18038, A2 => n16621, B1 => n16864, B2 => 
                           n16622, ZN => n4262);
   U15180 : OAI22_X1 port map( A1 => n18039, A2 => n16619, B1 => n16865, B2 => 
                           n16622, ZN => n4261);
   U15181 : OAI22_X1 port map( A1 => n18755, A2 => n16619, B1 => n16866, B2 => 
                           n16622, ZN => n4260);
   U15182 : OAI22_X1 port map( A1 => n18333, A2 => n16621, B1 => n16867, B2 => 
                           n16622, ZN => n4259);
   U15183 : OAI22_X1 port map( A1 => n18334, A2 => n16619, B1 => n16868, B2 => 
                           n16622, ZN => n4258);
   U15184 : OAI22_X1 port map( A1 => n18040, A2 => n16621, B1 => n16869, B2 => 
                           n16622, ZN => n4257);
   U15185 : OAI22_X1 port map( A1 => n18335, A2 => n16619, B1 => n16870, B2 => 
                           n16622, ZN => n4256);
   U15186 : OAI22_X1 port map( A1 => n18041, A2 => n16621, B1 => n16871, B2 => 
                           n16622, ZN => n4255);
   U15187 : OAI22_X1 port map( A1 => n18042, A2 => n16621, B1 => n16872, B2 => 
                           n16622, ZN => n4254);
   U15188 : OAI22_X1 port map( A1 => n18756, A2 => n16619, B1 => n16873, B2 => 
                           n16622, ZN => n4253);
   U15189 : OAI22_X1 port map( A1 => n18336, A2 => n16619, B1 => n16874, B2 => 
                           n16620, ZN => n4252);
   U15190 : OAI22_X1 port map( A1 => n18337, A2 => n16621, B1 => n16875, B2 => 
                           n16622, ZN => n4251);
   U15191 : OAI22_X1 port map( A1 => n18757, A2 => n16619, B1 => n16876, B2 => 
                           n16622, ZN => n4250);
   U15192 : OAI22_X1 port map( A1 => n18043, A2 => n16621, B1 => n16878, B2 => 
                           n16620, ZN => n4249);
   U15193 : OAI22_X1 port map( A1 => n18044, A2 => n16619, B1 => n16881, B2 => 
                           n16622, ZN => n4248);
   U15194 : INV_X1 port map( A => ADD_WR(2), ZN => n16638);
   U15195 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n16638, 
                           ZN => n16734);
   U15196 : NAND2_X1 port map( A1 => n16639, A2 => n16734, ZN => n16625);
   U15197 : NAND2_X1 port map( A1 => n13731, A2 => n16624, ZN => n16626);
   U15198 : CLKBUF_X2 port map( A => n16625, Z => n16624);
   U15199 : OAI22_X1 port map( A1 => n16885, A2 => n16626, B1 => n16815, B2 => 
                           n16624, ZN => n4247);
   U15200 : CLKBUF_X2 port map( A => n16626, Z => n16623);
   U15201 : OAI22_X1 port map( A1 => n18338, A2 => n16623, B1 => n16746, B2 => 
                           n16625, ZN => n4246);
   U15202 : OAI22_X1 port map( A1 => n18045, A2 => n16626, B1 => n16747, B2 => 
                           n16625, ZN => n4245);
   U15203 : OAI22_X1 port map( A1 => n18339, A2 => n16623, B1 => n16748, B2 => 
                           n16624, ZN => n4244);
   U15204 : OAI22_X1 port map( A1 => n18046, A2 => n16623, B1 => n16749, B2 => 
                           n16625, ZN => n4243);
   U15205 : OAI22_X1 port map( A1 => n18340, A2 => n16623, B1 => n16750, B2 => 
                           n16624, ZN => n4242);
   U15206 : OAI22_X1 port map( A1 => n18341, A2 => n16623, B1 => n16751, B2 => 
                           n16625, ZN => n4241);
   U15207 : OAI22_X1 port map( A1 => n18047, A2 => n16623, B1 => n16752, B2 => 
                           n16625, ZN => n4240);
   U15208 : OAI22_X1 port map( A1 => n18048, A2 => n16623, B1 => n16753, B2 => 
                           n16624, ZN => n4239);
   U15209 : OAI22_X1 port map( A1 => n18342, A2 => n16623, B1 => n16754, B2 => 
                           n16625, ZN => n4238);
   U15210 : OAI22_X1 port map( A1 => n18343, A2 => n16623, B1 => n16755, B2 => 
                           n16624, ZN => n4237);
   U15211 : OAI22_X1 port map( A1 => n18049, A2 => n16623, B1 => n16756, B2 => 
                           n16624, ZN => n4236);
   U15212 : OAI22_X1 port map( A1 => n18050, A2 => n16626, B1 => n16757, B2 => 
                           n16625, ZN => n4235);
   U15213 : OAI22_X1 port map( A1 => n18051, A2 => n16623, B1 => n16758, B2 => 
                           n16624, ZN => n4234);
   U15214 : OAI22_X1 port map( A1 => n18052, A2 => n16623, B1 => n16759, B2 => 
                           n16625, ZN => n4233);
   U15215 : OAI22_X1 port map( A1 => n18053, A2 => n16626, B1 => n16760, B2 => 
                           n16624, ZN => n4232);
   U15216 : OAI22_X1 port map( A1 => n18758, A2 => n16626, B1 => n16761, B2 => 
                           n16625, ZN => n4231);
   U15217 : OAI22_X1 port map( A1 => n18054, A2 => n16623, B1 => n16762, B2 => 
                           n16624, ZN => n4230);
   U15218 : OAI22_X1 port map( A1 => n18055, A2 => n16623, B1 => n16763, B2 => 
                           n16625, ZN => n4229);
   U15219 : OAI22_X1 port map( A1 => n18344, A2 => n16626, B1 => n16764, B2 => 
                           n16624, ZN => n4228);
   U15220 : OAI22_X1 port map( A1 => n18056, A2 => n16626, B1 => n16765, B2 => 
                           n16625, ZN => n4227);
   U15221 : OAI22_X1 port map( A1 => n18057, A2 => n16623, B1 => n16766, B2 => 
                           n16624, ZN => n4226);
   U15222 : OAI22_X1 port map( A1 => n18345, A2 => n16623, B1 => n16767, B2 => 
                           n16624, ZN => n4225);
   U15223 : OAI22_X1 port map( A1 => n18058, A2 => n16623, B1 => n16768, B2 => 
                           n16625, ZN => n4224);
   U15224 : OAI22_X1 port map( A1 => n18346, A2 => n16623, B1 => n16769, B2 => 
                           n16624, ZN => n4223);
   U15225 : OAI22_X1 port map( A1 => n18347, A2 => n16626, B1 => n16770, B2 => 
                           n16625, ZN => n4222);
   U15226 : OAI22_X1 port map( A1 => n18348, A2 => n16623, B1 => n16771, B2 => 
                           n16625, ZN => n4221);
   U15227 : OAI22_X1 port map( A1 => n18059, A2 => n16626, B1 => n16772, B2 => 
                           n16625, ZN => n4220);
   U15228 : OAI22_X1 port map( A1 => n18349, A2 => n16623, B1 => n16773, B2 => 
                           n16625, ZN => n4219);
   U15229 : OAI22_X1 port map( A1 => n18060, A2 => n16626, B1 => n16774, B2 => 
                           n16625, ZN => n4218);
   U15230 : OAI22_X1 port map( A1 => n18350, A2 => n16623, B1 => n16775, B2 => 
                           n16625, ZN => n4217);
   U15231 : OAI22_X1 port map( A1 => n18351, A2 => n16626, B1 => n16776, B2 => 
                           n16625, ZN => n4216);
   U15232 : OAI22_X1 port map( A1 => n18759, A2 => n16623, B1 => n16777, B2 => 
                           n16625, ZN => n4215);
   U15233 : OAI22_X1 port map( A1 => n18352, A2 => n16626, B1 => n16778, B2 => 
                           n16625, ZN => n4214);
   U15234 : OAI22_X1 port map( A1 => n18061, A2 => n16623, B1 => n16779, B2 => 
                           n16625, ZN => n4213);
   U15235 : OAI22_X1 port map( A1 => n18353, A2 => n16626, B1 => n16781, B2 => 
                           n16624, ZN => n4212);
   U15236 : OAI22_X1 port map( A1 => n17194, A2 => n16626, B1 => n16782, B2 => 
                           n16624, ZN => n4211);
   U15237 : OAI22_X1 port map( A1 => n17810, A2 => n16623, B1 => n16783, B2 => 
                           n16624, ZN => n4210);
   U15238 : OAI22_X1 port map( A1 => n17422, A2 => n16626, B1 => n16784, B2 => 
                           n16624, ZN => n4209);
   U15239 : OAI22_X1 port map( A1 => n17423, A2 => n16623, B1 => n16785, B2 => 
                           n16624, ZN => n4208);
   U15240 : OAI22_X1 port map( A1 => n17424, A2 => n16626, B1 => n16786, B2 => 
                           n16624, ZN => n4207);
   U15241 : OAI22_X1 port map( A1 => n17195, A2 => n16623, B1 => n16787, B2 => 
                           n16624, ZN => n4206);
   U15242 : OAI22_X1 port map( A1 => n17425, A2 => n16623, B1 => n16788, B2 => 
                           n16624, ZN => n4205);
   U15243 : OAI22_X1 port map( A1 => n17811, A2 => n16623, B1 => n16789, B2 => 
                           n16624, ZN => n4204);
   U15244 : OAI22_X1 port map( A1 => n17426, A2 => n16623, B1 => n16790, B2 => 
                           n16624, ZN => n4203);
   U15245 : OAI22_X1 port map( A1 => n17196, A2 => n16623, B1 => n16791, B2 => 
                           n16624, ZN => n4202);
   U15246 : OAI22_X1 port map( A1 => n17812, A2 => n16623, B1 => n16792, B2 => 
                           n16624, ZN => n4201);
   U15247 : OAI22_X1 port map( A1 => n17197, A2 => n16623, B1 => n16793, B2 => 
                           n16624, ZN => n4200);
   U15248 : OAI22_X1 port map( A1 => n18354, A2 => n16626, B1 => n16794, B2 => 
                           n16624, ZN => n4199);
   U15249 : OAI22_X1 port map( A1 => n18355, A2 => n16626, B1 => n16795, B2 => 
                           n16624, ZN => n4198);
   U15250 : OAI22_X1 port map( A1 => n18062, A2 => n16623, B1 => n16796, B2 => 
                           n16624, ZN => n4197);
   U15251 : OAI22_X1 port map( A1 => n18356, A2 => n16623, B1 => n16797, B2 => 
                           n16624, ZN => n4196);
   U15252 : OAI22_X1 port map( A1 => n18357, A2 => n16626, B1 => n16798, B2 => 
                           n16624, ZN => n4195);
   U15253 : OAI22_X1 port map( A1 => n18358, A2 => n16623, B1 => n16799, B2 => 
                           n16624, ZN => n4194);
   U15254 : OAI22_X1 port map( A1 => n18359, A2 => n16626, B1 => n16800, B2 => 
                           n16624, ZN => n4193);
   U15255 : OAI22_X1 port map( A1 => n18360, A2 => n16623, B1 => n16801, B2 => 
                           n16624, ZN => n4192);
   U15256 : OAI22_X1 port map( A1 => n18760, A2 => n16626, B1 => n16802, B2 => 
                           n16624, ZN => n4191);
   U15257 : OAI22_X1 port map( A1 => n18761, A2 => n16626, B1 => n16803, B2 => 
                           n16624, ZN => n4190);
   U15258 : OAI22_X1 port map( A1 => n18063, A2 => n16623, B1 => n16804, B2 => 
                           n16624, ZN => n4189);
   U15259 : OAI22_X1 port map( A1 => n18064, A2 => n16623, B1 => n16805, B2 => 
                           n16625, ZN => n4188);
   U15260 : OAI22_X1 port map( A1 => n18762, A2 => n16626, B1 => n16806, B2 => 
                           n16624, ZN => n4187);
   U15261 : OAI22_X1 port map( A1 => n18361, A2 => n16623, B1 => n16808, B2 => 
                           n16624, ZN => n4186);
   U15262 : OAI22_X1 port map( A1 => n18362, A2 => n16626, B1 => n16810, B2 => 
                           n16625, ZN => n4185);
   U15263 : OAI22_X1 port map( A1 => n18363, A2 => n16623, B1 => n16812, B2 => 
                           n16624, ZN => n4184);
   U15264 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => n16627, A3 => n16638, ZN 
                           => n16739);
   U15265 : NAND2_X1 port map( A1 => n16639, A2 => n16739, ZN => n16629);
   U15266 : CLKBUF_X2 port map( A => n16629, Z => n16631);
   U15267 : NAND2_X1 port map( A1 => n13731, A2 => n16631, ZN => n16630);
   U15268 : OAI22_X1 port map( A1 => n16886, A2 => n16630, B1 => n16745, B2 => 
                           n16631, ZN => n4183);
   U15269 : CLKBUF_X2 port map( A => n16630, Z => n16628);
   U15270 : OAI22_X1 port map( A1 => n18364, A2 => n16628, B1 => n16816, B2 => 
                           n16629, ZN => n4182);
   U15271 : OAI22_X1 port map( A1 => n18365, A2 => n16630, B1 => n16817, B2 => 
                           n16631, ZN => n4181);
   U15272 : OAI22_X1 port map( A1 => n18366, A2 => n16628, B1 => n16818, B2 => 
                           n16629, ZN => n4180);
   U15273 : OAI22_X1 port map( A1 => n18367, A2 => n16628, B1 => n16819, B2 => 
                           n16629, ZN => n4179);
   U15274 : OAI22_X1 port map( A1 => n18763, A2 => n16628, B1 => n16820, B2 => 
                           n16631, ZN => n4178);
   U15275 : OAI22_X1 port map( A1 => n18368, A2 => n16628, B1 => n16821, B2 => 
                           n16629, ZN => n4177);
   U15276 : OAI22_X1 port map( A1 => n18764, A2 => n16628, B1 => n16822, B2 => 
                           n16631, ZN => n4176);
   U15277 : OAI22_X1 port map( A1 => n18765, A2 => n16628, B1 => n16823, B2 => 
                           n16631, ZN => n4175);
   U15278 : OAI22_X1 port map( A1 => n18766, A2 => n16628, B1 => n16824, B2 => 
                           n16631, ZN => n4174);
   U15279 : OAI22_X1 port map( A1 => n18369, A2 => n16628, B1 => n16825, B2 => 
                           n16631, ZN => n4173);
   U15280 : OAI22_X1 port map( A1 => n18767, A2 => n16628, B1 => n16826, B2 => 
                           n16631, ZN => n4172);
   U15281 : OAI22_X1 port map( A1 => n18065, A2 => n16630, B1 => n16827, B2 => 
                           n16629, ZN => n4171);
   U15282 : OAI22_X1 port map( A1 => n18768, A2 => n16628, B1 => n16828, B2 => 
                           n16629, ZN => n4170);
   U15283 : OAI22_X1 port map( A1 => n18370, A2 => n16628, B1 => n16829, B2 => 
                           n16629, ZN => n4169);
   U15284 : OAI22_X1 port map( A1 => n18371, A2 => n16630, B1 => n16830, B2 => 
                           n16631, ZN => n4168);
   U15285 : OAI22_X1 port map( A1 => n18769, A2 => n16630, B1 => n16831, B2 => 
                           n16629, ZN => n4167);
   U15286 : OAI22_X1 port map( A1 => n18770, A2 => n16628, B1 => n16832, B2 => 
                           n16629, ZN => n4166);
   U15287 : OAI22_X1 port map( A1 => n18372, A2 => n16628, B1 => n16833, B2 => 
                           n16629, ZN => n4165);
   U15288 : OAI22_X1 port map( A1 => n18373, A2 => n16630, B1 => n16834, B2 => 
                           n16631, ZN => n4164);
   U15289 : OAI22_X1 port map( A1 => n18374, A2 => n16630, B1 => n16835, B2 => 
                           n16629, ZN => n4163);
   U15290 : OAI22_X1 port map( A1 => n18771, A2 => n16628, B1 => n16836, B2 => 
                           n16631, ZN => n4162);
   U15291 : OAI22_X1 port map( A1 => n18772, A2 => n16628, B1 => n16837, B2 => 
                           n16631, ZN => n4161);
   U15292 : OAI22_X1 port map( A1 => n18773, A2 => n16628, B1 => n16838, B2 => 
                           n16629, ZN => n4160);
   U15293 : OAI22_X1 port map( A1 => n18774, A2 => n16628, B1 => n16839, B2 => 
                           n16631, ZN => n4159);
   U15294 : OAI22_X1 port map( A1 => n18775, A2 => n16630, B1 => n16840, B2 => 
                           n16629, ZN => n4158);
   U15295 : OAI22_X1 port map( A1 => n18375, A2 => n16628, B1 => n16841, B2 => 
                           n16629, ZN => n4157);
   U15296 : OAI22_X1 port map( A1 => n18776, A2 => n16630, B1 => n16842, B2 => 
                           n16629, ZN => n4156);
   U15297 : OAI22_X1 port map( A1 => n18777, A2 => n16628, B1 => n16843, B2 => 
                           n16629, ZN => n4155);
   U15298 : OAI22_X1 port map( A1 => n18376, A2 => n16630, B1 => n16844, B2 => 
                           n16629, ZN => n4154);
   U15299 : OAI22_X1 port map( A1 => n18778, A2 => n16628, B1 => n16845, B2 => 
                           n16629, ZN => n4153);
   U15300 : OAI22_X1 port map( A1 => n18779, A2 => n16630, B1 => n16846, B2 => 
                           n16629, ZN => n4152);
   U15301 : OAI22_X1 port map( A1 => n18780, A2 => n16628, B1 => n16847, B2 => 
                           n16629, ZN => n4151);
   U15302 : OAI22_X1 port map( A1 => n18377, A2 => n16630, B1 => n16848, B2 => 
                           n16629, ZN => n4150);
   U15303 : OAI22_X1 port map( A1 => n18378, A2 => n16628, B1 => n16849, B2 => 
                           n16629, ZN => n4149);
   U15304 : OAI22_X1 port map( A1 => n18379, A2 => n16630, B1 => n16850, B2 => 
                           n16631, ZN => n4148);
   U15305 : OAI22_X1 port map( A1 => n17427, A2 => n16630, B1 => n16851, B2 => 
                           n16631, ZN => n4147);
   U15306 : OAI22_X1 port map( A1 => n17428, A2 => n16628, B1 => n16852, B2 => 
                           n16631, ZN => n4146);
   U15307 : OAI22_X1 port map( A1 => n17429, A2 => n16630, B1 => n16853, B2 => 
                           n16631, ZN => n4145);
   U15308 : OAI22_X1 port map( A1 => n17430, A2 => n16628, B1 => n16854, B2 => 
                           n16631, ZN => n4144);
   U15309 : OAI22_X1 port map( A1 => n17198, A2 => n16630, B1 => n16855, B2 => 
                           n16631, ZN => n4143);
   U15310 : OAI22_X1 port map( A1 => n17813, A2 => n16628, B1 => n16856, B2 => 
                           n16631, ZN => n4142);
   U15311 : OAI22_X1 port map( A1 => n17814, A2 => n16628, B1 => n16857, B2 => 
                           n16631, ZN => n4141);
   U15312 : OAI22_X1 port map( A1 => n17815, A2 => n16628, B1 => n16858, B2 => 
                           n16631, ZN => n4140);
   U15313 : OAI22_X1 port map( A1 => n17816, A2 => n16628, B1 => n16859, B2 => 
                           n16631, ZN => n4139);
   U15314 : OAI22_X1 port map( A1 => n17431, A2 => n16628, B1 => n16860, B2 => 
                           n16631, ZN => n4138);
   U15315 : OAI22_X1 port map( A1 => n17199, A2 => n16628, B1 => n16861, B2 => 
                           n16631, ZN => n4137);
   U15316 : OAI22_X1 port map( A1 => n17817, A2 => n16628, B1 => n16862, B2 => 
                           n16631, ZN => n4136);
   U15317 : OAI22_X1 port map( A1 => n18066, A2 => n16630, B1 => n16863, B2 => 
                           n16631, ZN => n4135);
   U15318 : OAI22_X1 port map( A1 => n18781, A2 => n16630, B1 => n16864, B2 => 
                           n16631, ZN => n4134);
   U15319 : OAI22_X1 port map( A1 => n18067, A2 => n16628, B1 => n16865, B2 => 
                           n16631, ZN => n4133);
   U15320 : OAI22_X1 port map( A1 => n18380, A2 => n16628, B1 => n16866, B2 => 
                           n16631, ZN => n4132);
   U15321 : OAI22_X1 port map( A1 => n18068, A2 => n16630, B1 => n16867, B2 => 
                           n16631, ZN => n4131);
   U15322 : OAI22_X1 port map( A1 => n18782, A2 => n16628, B1 => n16868, B2 => 
                           n16631, ZN => n4130);
   U15323 : OAI22_X1 port map( A1 => n18783, A2 => n16630, B1 => n16869, B2 => 
                           n16631, ZN => n4129);
   U15324 : OAI22_X1 port map( A1 => n18784, A2 => n16628, B1 => n16870, B2 => 
                           n16631, ZN => n4128);
   U15325 : OAI22_X1 port map( A1 => n18069, A2 => n16630, B1 => n16871, B2 => 
                           n16631, ZN => n4127);
   U15326 : OAI22_X1 port map( A1 => n18381, A2 => n16630, B1 => n16872, B2 => 
                           n16631, ZN => n4126);
   U15327 : OAI22_X1 port map( A1 => n18382, A2 => n16628, B1 => n16873, B2 => 
                           n16631, ZN => n4125);
   U15328 : OAI22_X1 port map( A1 => n18383, A2 => n16628, B1 => n16874, B2 => 
                           n16629, ZN => n4124);
   U15329 : OAI22_X1 port map( A1 => n18384, A2 => n16630, B1 => n16875, B2 => 
                           n16631, ZN => n4123);
   U15330 : OAI22_X1 port map( A1 => n18385, A2 => n16628, B1 => n16876, B2 => 
                           n16631, ZN => n4122);
   U15331 : OAI22_X1 port map( A1 => n18386, A2 => n16630, B1 => n16878, B2 => 
                           n16629, ZN => n4121);
   U15332 : OAI22_X1 port map( A1 => n18387, A2 => n16628, B1 => n16881, B2 => 
                           n16631, ZN => n4120);
   U15333 : NOR2_X1 port map( A1 => n16638, A2 => n16632, ZN => n16744);
   U15334 : NAND2_X1 port map( A1 => n16639, A2 => n16744, ZN => n16634);
   U15335 : CLKBUF_X2 port map( A => n16634, Z => n16636);
   U15336 : NAND2_X1 port map( A1 => n13731, A2 => n16636, ZN => n16635);
   U15337 : OAI22_X1 port map( A1 => n16964, A2 => n16635, B1 => n16815, B2 => 
                           n16636, ZN => n4119);
   U15338 : CLKBUF_X2 port map( A => n16635, Z => n16633);
   U15339 : OAI22_X1 port map( A1 => n18388, A2 => n16633, B1 => n16746, B2 => 
                           n16634, ZN => n4118);
   U15340 : OAI22_X1 port map( A1 => n18785, A2 => n16635, B1 => n16747, B2 => 
                           n16636, ZN => n4117);
   U15341 : OAI22_X1 port map( A1 => n18389, A2 => n16633, B1 => n16748, B2 => 
                           n16634, ZN => n4116);
   U15342 : OAI22_X1 port map( A1 => n18390, A2 => n16633, B1 => n16749, B2 => 
                           n16634, ZN => n4115);
   U15343 : OAI22_X1 port map( A1 => n18391, A2 => n16633, B1 => n16750, B2 => 
                           n16636, ZN => n4114);
   U15344 : OAI22_X1 port map( A1 => n18392, A2 => n16633, B1 => n16751, B2 => 
                           n16634, ZN => n4113);
   U15345 : OAI22_X1 port map( A1 => n18786, A2 => n16633, B1 => n16752, B2 => 
                           n16636, ZN => n4112);
   U15346 : OAI22_X1 port map( A1 => n18393, A2 => n16633, B1 => n16753, B2 => 
                           n16636, ZN => n4111);
   U15347 : OAI22_X1 port map( A1 => n18070, A2 => n16633, B1 => n16754, B2 => 
                           n16636, ZN => n4110);
   U15348 : OAI22_X1 port map( A1 => n18394, A2 => n16633, B1 => n16755, B2 => 
                           n16636, ZN => n4109);
   U15349 : OAI22_X1 port map( A1 => n18071, A2 => n16633, B1 => n16756, B2 => 
                           n16636, ZN => n4108);
   U15350 : OAI22_X1 port map( A1 => n18395, A2 => n16635, B1 => n16757, B2 => 
                           n16634, ZN => n4107);
   U15351 : OAI22_X1 port map( A1 => n18396, A2 => n16633, B1 => n16758, B2 => 
                           n16634, ZN => n4106);
   U15352 : OAI22_X1 port map( A1 => n18787, A2 => n16633, B1 => n16759, B2 => 
                           n16634, ZN => n4105);
   U15353 : OAI22_X1 port map( A1 => n18788, A2 => n16635, B1 => n16760, B2 => 
                           n16636, ZN => n4104);
   U15354 : OAI22_X1 port map( A1 => n18072, A2 => n16635, B1 => n16761, B2 => 
                           n16634, ZN => n4103);
   U15355 : OAI22_X1 port map( A1 => n18397, A2 => n16633, B1 => n16762, B2 => 
                           n16634, ZN => n4102);
   U15356 : OAI22_X1 port map( A1 => n18398, A2 => n16633, B1 => n16763, B2 => 
                           n16634, ZN => n4101);
   U15357 : OAI22_X1 port map( A1 => n18073, A2 => n16635, B1 => n16764, B2 => 
                           n16636, ZN => n4100);
   U15358 : OAI22_X1 port map( A1 => n18789, A2 => n16635, B1 => n16765, B2 => 
                           n16634, ZN => n4099);
   U15359 : OAI22_X1 port map( A1 => n18399, A2 => n16633, B1 => n16766, B2 => 
                           n16636, ZN => n4098);
   U15360 : OAI22_X1 port map( A1 => n18400, A2 => n16633, B1 => n16767, B2 => 
                           n16636, ZN => n4097);
   U15361 : OAI22_X1 port map( A1 => n18790, A2 => n16633, B1 => n16768, B2 => 
                           n16634, ZN => n4096);
   U15362 : OAI22_X1 port map( A1 => n18074, A2 => n16633, B1 => n16769, B2 => 
                           n16636, ZN => n4095);
   U15363 : OAI22_X1 port map( A1 => n18075, A2 => n16635, B1 => n16770, B2 => 
                           n16634, ZN => n4094);
   U15364 : OAI22_X1 port map( A1 => n18791, A2 => n16633, B1 => n16771, B2 => 
                           n16634, ZN => n4093);
   U15365 : OAI22_X1 port map( A1 => n18076, A2 => n16635, B1 => n16772, B2 => 
                           n16634, ZN => n4092);
   U15366 : OAI22_X1 port map( A1 => n18077, A2 => n16633, B1 => n16773, B2 => 
                           n16634, ZN => n4091);
   U15367 : OAI22_X1 port map( A1 => n18401, A2 => n16635, B1 => n16774, B2 => 
                           n16634, ZN => n4090);
   U15368 : OAI22_X1 port map( A1 => n18402, A2 => n16633, B1 => n16775, B2 => 
                           n16634, ZN => n4089);
   U15369 : OAI22_X1 port map( A1 => n18078, A2 => n16635, B1 => n16776, B2 => 
                           n16634, ZN => n4088);
   U15370 : OAI22_X1 port map( A1 => n18079, A2 => n16633, B1 => n16777, B2 => 
                           n16634, ZN => n4087);
   U15371 : OAI22_X1 port map( A1 => n18403, A2 => n16635, B1 => n16778, B2 => 
                           n16634, ZN => n4086);
   U15372 : OAI22_X1 port map( A1 => n18404, A2 => n16633, B1 => n16779, B2 => 
                           n16634, ZN => n4085);
   U15373 : OAI22_X1 port map( A1 => n18405, A2 => n16635, B1 => n16781, B2 => 
                           n16636, ZN => n4084);
   U15374 : OAI22_X1 port map( A1 => n17432, A2 => n16635, B1 => n16782, B2 => 
                           n16636, ZN => n4083);
   U15375 : OAI22_X1 port map( A1 => n17200, A2 => n16633, B1 => n16783, B2 => 
                           n16636, ZN => n4082);
   U15376 : OAI22_X1 port map( A1 => n17818, A2 => n16635, B1 => n16784, B2 => 
                           n16636, ZN => n4081);
   U15377 : OAI22_X1 port map( A1 => n17433, A2 => n16633, B1 => n16785, B2 => 
                           n16636, ZN => n4080);
   U15378 : OAI22_X1 port map( A1 => n17819, A2 => n16635, B1 => n16786, B2 => 
                           n16636, ZN => n4079);
   U15379 : OAI22_X1 port map( A1 => n17434, A2 => n16633, B1 => n16787, B2 => 
                           n16636, ZN => n4078);
   U15380 : OAI22_X1 port map( A1 => n17435, A2 => n16633, B1 => n16788, B2 => 
                           n16636, ZN => n4077);
   U15381 : OAI22_X1 port map( A1 => n17436, A2 => n16633, B1 => n16789, B2 => 
                           n16636, ZN => n4076);
   U15382 : OAI22_X1 port map( A1 => n17201, A2 => n16633, B1 => n16790, B2 => 
                           n16636, ZN => n4075);
   U15383 : OAI22_X1 port map( A1 => n17437, A2 => n16633, B1 => n16791, B2 => 
                           n16636, ZN => n4074);
   U15384 : OAI22_X1 port map( A1 => n17202, A2 => n16633, B1 => n16792, B2 => 
                           n16636, ZN => n4073);
   U15385 : OAI22_X1 port map( A1 => n17203, A2 => n16633, B1 => n16793, B2 => 
                           n16636, ZN => n4072);
   U15386 : OAI22_X1 port map( A1 => n18406, A2 => n16635, B1 => n16794, B2 => 
                           n16636, ZN => n4071);
   U15387 : OAI22_X1 port map( A1 => n18407, A2 => n16635, B1 => n16795, B2 => 
                           n16636, ZN => n4070);
   U15388 : OAI22_X1 port map( A1 => n18792, A2 => n16633, B1 => n16796, B2 => 
                           n16636, ZN => n4069);
   U15389 : OAI22_X1 port map( A1 => n18408, A2 => n16633, B1 => n16797, B2 => 
                           n16636, ZN => n4068);
   U15390 : OAI22_X1 port map( A1 => n18409, A2 => n16635, B1 => n16798, B2 => 
                           n16636, ZN => n4067);
   U15391 : OAI22_X1 port map( A1 => n18410, A2 => n16633, B1 => n16799, B2 => 
                           n16636, ZN => n4066);
   U15392 : OAI22_X1 port map( A1 => n18411, A2 => n16635, B1 => n16800, B2 => 
                           n16636, ZN => n4065);
   U15393 : OAI22_X1 port map( A1 => n18080, A2 => n16633, B1 => n16801, B2 => 
                           n16636, ZN => n4064);
   U15394 : OAI22_X1 port map( A1 => n18793, A2 => n16635, B1 => n16802, B2 => 
                           n16636, ZN => n4063);
   U15395 : OAI22_X1 port map( A1 => n18412, A2 => n16635, B1 => n16803, B2 => 
                           n16636, ZN => n4062);
   U15396 : OAI22_X1 port map( A1 => n18413, A2 => n16633, B1 => n16804, B2 => 
                           n16636, ZN => n4061);
   U15397 : OAI22_X1 port map( A1 => n18414, A2 => n16633, B1 => n16805, B2 => 
                           n16634, ZN => n4060);
   U15398 : OAI22_X1 port map( A1 => n18081, A2 => n16635, B1 => n16806, B2 => 
                           n16636, ZN => n4059);
   U15399 : OAI22_X1 port map( A1 => n18415, A2 => n16633, B1 => n16808, B2 => 
                           n16636, ZN => n4058);
   U15400 : OAI22_X1 port map( A1 => n18794, A2 => n16635, B1 => n16810, B2 => 
                           n16634, ZN => n4057);
   U15401 : OAI22_X1 port map( A1 => n18795, A2 => n16633, B1 => n16812, B2 => 
                           n16636, ZN => n4056);
   U15402 : NOR2_X1 port map( A1 => n16638, A2 => n16637, ZN => n16814);
   U15403 : NAND2_X1 port map( A1 => n16639, A2 => n16814, ZN => n16641);
   U15404 : CLKBUF_X2 port map( A => n16641, Z => n16643);
   U15405 : NAND2_X1 port map( A1 => n13731, A2 => n16643, ZN => n16642);
   U15406 : OAI22_X1 port map( A1 => n17107, A2 => n16642, B1 => n16745, B2 => 
                           n16643, ZN => n4055);
   U15407 : CLKBUF_X2 port map( A => n16642, Z => n16640);
   U15408 : OAI22_X1 port map( A1 => n18416, A2 => n16640, B1 => n16816, B2 => 
                           n16641, ZN => n4054);
   U15409 : OAI22_X1 port map( A1 => n18417, A2 => n16642, B1 => n16817, B2 => 
                           n16643, ZN => n4053);
   U15410 : OAI22_X1 port map( A1 => n18418, A2 => n16640, B1 => n16818, B2 => 
                           n16641, ZN => n4052);
   U15411 : OAI22_X1 port map( A1 => n18082, A2 => n16640, B1 => n16819, B2 => 
                           n16641, ZN => n4051);
   U15412 : OAI22_X1 port map( A1 => n18083, A2 => n16640, B1 => n16820, B2 => 
                           n16643, ZN => n4050);
   U15413 : OAI22_X1 port map( A1 => n18419, A2 => n16640, B1 => n16821, B2 => 
                           n16641, ZN => n4049);
   U15414 : OAI22_X1 port map( A1 => n18420, A2 => n16640, B1 => n16822, B2 => 
                           n16643, ZN => n4048);
   U15415 : OAI22_X1 port map( A1 => n18421, A2 => n16640, B1 => n16823, B2 => 
                           n16643, ZN => n4047);
   U15416 : OAI22_X1 port map( A1 => n18084, A2 => n16640, B1 => n16824, B2 => 
                           n16643, ZN => n4046);
   U15417 : OAI22_X1 port map( A1 => n18085, A2 => n16640, B1 => n16825, B2 => 
                           n16643, ZN => n4045);
   U15418 : OAI22_X1 port map( A1 => n18422, A2 => n16640, B1 => n16826, B2 => 
                           n16643, ZN => n4044);
   U15419 : OAI22_X1 port map( A1 => n18796, A2 => n16642, B1 => n16827, B2 => 
                           n16641, ZN => n4043);
   U15420 : OAI22_X1 port map( A1 => n18086, A2 => n16640, B1 => n16828, B2 => 
                           n16641, ZN => n4042);
   U15421 : OAI22_X1 port map( A1 => n18423, A2 => n16640, B1 => n16829, B2 => 
                           n16641, ZN => n4041);
   U15422 : OAI22_X1 port map( A1 => n18087, A2 => n16642, B1 => n16830, B2 => 
                           n16643, ZN => n4040);
   U15423 : OAI22_X1 port map( A1 => n18088, A2 => n16642, B1 => n16831, B2 => 
                           n16641, ZN => n4039);
   U15424 : OAI22_X1 port map( A1 => n18424, A2 => n16640, B1 => n16832, B2 => 
                           n16641, ZN => n4038);
   U15425 : OAI22_X1 port map( A1 => n18089, A2 => n16640, B1 => n16833, B2 => 
                           n16641, ZN => n4037);
   U15426 : OAI22_X1 port map( A1 => n18797, A2 => n16642, B1 => n16834, B2 => 
                           n16643, ZN => n4036);
   U15427 : OAI22_X1 port map( A1 => n18090, A2 => n16642, B1 => n16835, B2 => 
                           n16641, ZN => n4035);
   U15428 : OAI22_X1 port map( A1 => n18425, A2 => n16640, B1 => n16836, B2 => 
                           n16643, ZN => n4034);
   U15429 : OAI22_X1 port map( A1 => n18426, A2 => n16640, B1 => n16837, B2 => 
                           n16643, ZN => n4033);
   U15430 : OAI22_X1 port map( A1 => n18427, A2 => n16640, B1 => n16838, B2 => 
                           n16641, ZN => n4032);
   U15431 : OAI22_X1 port map( A1 => n18428, A2 => n16640, B1 => n16839, B2 => 
                           n16643, ZN => n4031);
   U15432 : OAI22_X1 port map( A1 => n18091, A2 => n16642, B1 => n16840, B2 => 
                           n16641, ZN => n4030);
   U15433 : OAI22_X1 port map( A1 => n18092, A2 => n16640, B1 => n16841, B2 => 
                           n16641, ZN => n4029);
   U15434 : OAI22_X1 port map( A1 => n18429, A2 => n16642, B1 => n16842, B2 => 
                           n16641, ZN => n4028);
   U15435 : OAI22_X1 port map( A1 => n18093, A2 => n16640, B1 => n16843, B2 => 
                           n16641, ZN => n4027);
   U15436 : OAI22_X1 port map( A1 => n18430, A2 => n16642, B1 => n16844, B2 => 
                           n16641, ZN => n4026);
   U15437 : OAI22_X1 port map( A1 => n18431, A2 => n16640, B1 => n16845, B2 => 
                           n16641, ZN => n4025);
   U15438 : OAI22_X1 port map( A1 => n18432, A2 => n16642, B1 => n16846, B2 => 
                           n16641, ZN => n4024);
   U15439 : OAI22_X1 port map( A1 => n18433, A2 => n16640, B1 => n16847, B2 => 
                           n16641, ZN => n4023);
   U15440 : OAI22_X1 port map( A1 => n18094, A2 => n16642, B1 => n16848, B2 => 
                           n16641, ZN => n4022);
   U15441 : OAI22_X1 port map( A1 => n18434, A2 => n16640, B1 => n16849, B2 => 
                           n16641, ZN => n4021);
   U15442 : OAI22_X1 port map( A1 => n18095, A2 => n16642, B1 => n16850, B2 => 
                           n16643, ZN => n4020);
   U15443 : OAI22_X1 port map( A1 => n17438, A2 => n16642, B1 => n16851, B2 => 
                           n16643, ZN => n4019);
   U15444 : OAI22_X1 port map( A1 => n17204, A2 => n16640, B1 => n16852, B2 => 
                           n16643, ZN => n4018);
   U15445 : OAI22_X1 port map( A1 => n17205, A2 => n16642, B1 => n16853, B2 => 
                           n16643, ZN => n4017);
   U15446 : OAI22_X1 port map( A1 => n17206, A2 => n16640, B1 => n16854, B2 => 
                           n16643, ZN => n4016);
   U15447 : OAI22_X1 port map( A1 => n17207, A2 => n16642, B1 => n16855, B2 => 
                           n16643, ZN => n4015);
   U15448 : OAI22_X1 port map( A1 => n17439, A2 => n16640, B1 => n16856, B2 => 
                           n16643, ZN => n4014);
   U15449 : OAI22_X1 port map( A1 => n17208, A2 => n16640, B1 => n16857, B2 => 
                           n16643, ZN => n4013);
   U15450 : OAI22_X1 port map( A1 => n17440, A2 => n16640, B1 => n16858, B2 => 
                           n16643, ZN => n4012);
   U15451 : OAI22_X1 port map( A1 => n17441, A2 => n16640, B1 => n16859, B2 => 
                           n16643, ZN => n4011);
   U15452 : OAI22_X1 port map( A1 => n17209, A2 => n16640, B1 => n16860, B2 => 
                           n16643, ZN => n4010);
   U15453 : OAI22_X1 port map( A1 => n17442, A2 => n16640, B1 => n16861, B2 => 
                           n16643, ZN => n4009);
   U15454 : OAI22_X1 port map( A1 => n17443, A2 => n16640, B1 => n16862, B2 => 
                           n16643, ZN => n4008);
   U15455 : OAI22_X1 port map( A1 => n18435, A2 => n16642, B1 => n16863, B2 => 
                           n16643, ZN => n4007);
   U15456 : OAI22_X1 port map( A1 => n18096, A2 => n16642, B1 => n16864, B2 => 
                           n16643, ZN => n4006);
   U15457 : OAI22_X1 port map( A1 => n18798, A2 => n16640, B1 => n16865, B2 => 
                           n16643, ZN => n4005);
   U15458 : OAI22_X1 port map( A1 => n18097, A2 => n16640, B1 => n16866, B2 => 
                           n16643, ZN => n4004);
   U15459 : OAI22_X1 port map( A1 => n18098, A2 => n16642, B1 => n16867, B2 => 
                           n16643, ZN => n4003);
   U15460 : OAI22_X1 port map( A1 => n18799, A2 => n16640, B1 => n16868, B2 => 
                           n16643, ZN => n4002);
   U15461 : OAI22_X1 port map( A1 => n18436, A2 => n16642, B1 => n16869, B2 => 
                           n16643, ZN => n4001);
   U15462 : OAI22_X1 port map( A1 => n18437, A2 => n16640, B1 => n16870, B2 => 
                           n16643, ZN => n4000);
   U15463 : OAI22_X1 port map( A1 => n18438, A2 => n16642, B1 => n16871, B2 => 
                           n16643, ZN => n3999);
   U15464 : OAI22_X1 port map( A1 => n18439, A2 => n16642, B1 => n16872, B2 => 
                           n16643, ZN => n3998);
   U15465 : OAI22_X1 port map( A1 => n18440, A2 => n16640, B1 => n16873, B2 => 
                           n16643, ZN => n3997);
   U15466 : OAI22_X1 port map( A1 => n18099, A2 => n16640, B1 => n16874, B2 => 
                           n16641, ZN => n3996);
   U15467 : OAI22_X1 port map( A1 => n18100, A2 => n16642, B1 => n16875, B2 => 
                           n16643, ZN => n3995);
   U15468 : OAI22_X1 port map( A1 => n18101, A2 => n16640, B1 => n16876, B2 => 
                           n16643, ZN => n3994);
   U15469 : OAI22_X1 port map( A1 => n18102, A2 => n16642, B1 => n16878, B2 => 
                           n16641, ZN => n3993);
   U15470 : OAI22_X1 port map( A1 => n18103, A2 => n16640, B1 => n16881, B2 => 
                           n16643, ZN => n3992);
   U15471 : NAND2_X1 port map( A1 => ENABLE, A2 => ADD_WR(3), ZN => n16713);
   U15472 : NOR2_X1 port map( A1 => n16644, A2 => n16713, ZN => n16673);
   U15473 : NAND2_X1 port map( A1 => n16714, A2 => n16673, ZN => n16646);
   U15474 : CLKBUF_X2 port map( A => n16646, Z => n16648);
   U15475 : NAND2_X1 port map( A1 => n13731, A2 => n16648, ZN => n16647);
   U15476 : OAI22_X1 port map( A1 => n16883, A2 => n16647, B1 => n16815, B2 => 
                           n16648, ZN => n3991);
   U15477 : CLKBUF_X2 port map( A => n16647, Z => n16645);
   U15478 : OAI22_X1 port map( A1 => n18441, A2 => n16645, B1 => n16816, B2 => 
                           n16646, ZN => n3990);
   U15479 : OAI22_X1 port map( A1 => n18442, A2 => n16647, B1 => n16817, B2 => 
                           n16648, ZN => n3989);
   U15480 : OAI22_X1 port map( A1 => n18800, A2 => n16645, B1 => n16818, B2 => 
                           n16646, ZN => n3988);
   U15481 : OAI22_X1 port map( A1 => n18104, A2 => n16645, B1 => n16819, B2 => 
                           n16646, ZN => n3987);
   U15482 : OAI22_X1 port map( A1 => n18443, A2 => n16645, B1 => n16820, B2 => 
                           n16648, ZN => n3986);
   U15483 : OAI22_X1 port map( A1 => n18444, A2 => n16645, B1 => n16821, B2 => 
                           n16646, ZN => n3985);
   U15484 : OAI22_X1 port map( A1 => n18445, A2 => n16645, B1 => n16822, B2 => 
                           n16648, ZN => n3984);
   U15485 : OAI22_X1 port map( A1 => n18105, A2 => n16645, B1 => n16823, B2 => 
                           n16648, ZN => n3983);
   U15486 : OAI22_X1 port map( A1 => n18446, A2 => n16645, B1 => n16824, B2 => 
                           n16648, ZN => n3982);
   U15487 : OAI22_X1 port map( A1 => n18447, A2 => n16645, B1 => n16825, B2 => 
                           n16648, ZN => n3981);
   U15488 : OAI22_X1 port map( A1 => n18106, A2 => n16645, B1 => n16826, B2 => 
                           n16648, ZN => n3980);
   U15489 : OAI22_X1 port map( A1 => n18448, A2 => n16647, B1 => n16827, B2 => 
                           n16646, ZN => n3979);
   U15490 : OAI22_X1 port map( A1 => n18449, A2 => n16645, B1 => n16828, B2 => 
                           n16646, ZN => n3978);
   U15491 : OAI22_X1 port map( A1 => n18450, A2 => n16645, B1 => n16829, B2 => 
                           n16646, ZN => n3977);
   U15492 : OAI22_X1 port map( A1 => n18451, A2 => n16647, B1 => n16830, B2 => 
                           n16648, ZN => n3976);
   U15493 : OAI22_X1 port map( A1 => n18452, A2 => n16647, B1 => n16831, B2 => 
                           n16646, ZN => n3975);
   U15494 : OAI22_X1 port map( A1 => n18453, A2 => n16645, B1 => n16832, B2 => 
                           n16646, ZN => n3974);
   U15495 : OAI22_X1 port map( A1 => n18454, A2 => n16645, B1 => n16833, B2 => 
                           n16646, ZN => n3973);
   U15496 : OAI22_X1 port map( A1 => n18801, A2 => n16647, B1 => n16834, B2 => 
                           n16648, ZN => n3972);
   U15497 : OAI22_X1 port map( A1 => n18107, A2 => n16647, B1 => n16835, B2 => 
                           n16646, ZN => n3971);
   U15498 : OAI22_X1 port map( A1 => n18802, A2 => n16645, B1 => n16836, B2 => 
                           n16648, ZN => n3970);
   U15499 : OAI22_X1 port map( A1 => n18455, A2 => n16645, B1 => n16837, B2 => 
                           n16648, ZN => n3969);
   U15500 : OAI22_X1 port map( A1 => n18108, A2 => n16645, B1 => n16838, B2 => 
                           n16646, ZN => n3968);
   U15501 : OAI22_X1 port map( A1 => n18456, A2 => n16645, B1 => n16839, B2 => 
                           n16648, ZN => n3967);
   U15502 : OAI22_X1 port map( A1 => n18457, A2 => n16647, B1 => n16840, B2 => 
                           n16646, ZN => n3966);
   U15503 : OAI22_X1 port map( A1 => n18109, A2 => n16645, B1 => n16841, B2 => 
                           n16646, ZN => n3965);
   U15504 : OAI22_X1 port map( A1 => n18458, A2 => n16647, B1 => n16842, B2 => 
                           n16646, ZN => n3964);
   U15505 : OAI22_X1 port map( A1 => n18110, A2 => n16645, B1 => n16843, B2 => 
                           n16646, ZN => n3963);
   U15506 : OAI22_X1 port map( A1 => n18459, A2 => n16647, B1 => n16844, B2 => 
                           n16646, ZN => n3962);
   U15507 : OAI22_X1 port map( A1 => n18111, A2 => n16645, B1 => n16845, B2 => 
                           n16646, ZN => n3961);
   U15508 : OAI22_X1 port map( A1 => n18112, A2 => n16647, B1 => n16846, B2 => 
                           n16646, ZN => n3960);
   U15509 : OAI22_X1 port map( A1 => n18113, A2 => n16645, B1 => n16847, B2 => 
                           n16646, ZN => n3959);
   U15510 : OAI22_X1 port map( A1 => n18460, A2 => n16647, B1 => n16848, B2 => 
                           n16646, ZN => n3958);
   U15511 : OAI22_X1 port map( A1 => n18461, A2 => n16645, B1 => n16849, B2 => 
                           n16646, ZN => n3957);
   U15512 : OAI22_X1 port map( A1 => n18114, A2 => n16647, B1 => n16850, B2 => 
                           n16648, ZN => n3956);
   U15513 : OAI22_X1 port map( A1 => n17820, A2 => n16647, B1 => n16851, B2 => 
                           n16648, ZN => n3955);
   U15514 : OAI22_X1 port map( A1 => n17821, A2 => n16645, B1 => n16852, B2 => 
                           n16648, ZN => n3954);
   U15515 : OAI22_X1 port map( A1 => n17444, A2 => n16647, B1 => n16853, B2 => 
                           n16648, ZN => n3953);
   U15516 : OAI22_X1 port map( A1 => n17445, A2 => n16645, B1 => n16854, B2 => 
                           n16648, ZN => n3952);
   U15517 : OAI22_X1 port map( A1 => n17446, A2 => n16647, B1 => n16855, B2 => 
                           n16648, ZN => n3951);
   U15518 : OAI22_X1 port map( A1 => n17447, A2 => n16645, B1 => n16856, B2 => 
                           n16648, ZN => n3950);
   U15519 : OAI22_X1 port map( A1 => n17210, A2 => n16645, B1 => n16857, B2 => 
                           n16648, ZN => n3949);
   U15520 : OAI22_X1 port map( A1 => n17448, A2 => n16645, B1 => n16858, B2 => 
                           n16648, ZN => n3948);
   U15521 : OAI22_X1 port map( A1 => n17211, A2 => n16645, B1 => n16859, B2 => 
                           n16648, ZN => n3947);
   U15522 : OAI22_X1 port map( A1 => n17822, A2 => n16645, B1 => n16860, B2 => 
                           n16648, ZN => n3946);
   U15523 : OAI22_X1 port map( A1 => n17449, A2 => n16645, B1 => n16861, B2 => 
                           n16648, ZN => n3945);
   U15524 : OAI22_X1 port map( A1 => n17450, A2 => n16645, B1 => n16862, B2 => 
                           n16648, ZN => n3944);
   U15525 : OAI22_X1 port map( A1 => n18462, A2 => n16647, B1 => n16863, B2 => 
                           n16648, ZN => n3943);
   U15526 : OAI22_X1 port map( A1 => n18803, A2 => n16647, B1 => n16864, B2 => 
                           n16648, ZN => n3942);
   U15527 : OAI22_X1 port map( A1 => n18115, A2 => n16645, B1 => n16865, B2 => 
                           n16648, ZN => n3941);
   U15528 : OAI22_X1 port map( A1 => n18463, A2 => n16645, B1 => n16866, B2 => 
                           n16648, ZN => n3940);
   U15529 : OAI22_X1 port map( A1 => n18464, A2 => n16647, B1 => n16867, B2 => 
                           n16648, ZN => n3939);
   U15530 : OAI22_X1 port map( A1 => n18116, A2 => n16645, B1 => n16868, B2 => 
                           n16648, ZN => n3938);
   U15531 : OAI22_X1 port map( A1 => n18465, A2 => n16647, B1 => n16869, B2 => 
                           n16648, ZN => n3937);
   U15532 : OAI22_X1 port map( A1 => n18466, A2 => n16645, B1 => n16870, B2 => 
                           n16648, ZN => n3936);
   U15533 : OAI22_X1 port map( A1 => n18117, A2 => n16647, B1 => n16871, B2 => 
                           n16648, ZN => n3935);
   U15534 : OAI22_X1 port map( A1 => n18467, A2 => n16647, B1 => n16872, B2 => 
                           n16648, ZN => n3934);
   U15535 : OAI22_X1 port map( A1 => n18468, A2 => n16645, B1 => n16873, B2 => 
                           n16648, ZN => n3933);
   U15536 : OAI22_X1 port map( A1 => n18118, A2 => n16645, B1 => n16874, B2 => 
                           n16646, ZN => n3932);
   U15537 : OAI22_X1 port map( A1 => n18469, A2 => n16647, B1 => n16875, B2 => 
                           n16648, ZN => n3931);
   U15538 : OAI22_X1 port map( A1 => n18119, A2 => n16645, B1 => n16876, B2 => 
                           n16648, ZN => n3930);
   U15539 : OAI22_X1 port map( A1 => n18470, A2 => n16647, B1 => n16878, B2 => 
                           n16646, ZN => n3929);
   U15540 : OAI22_X1 port map( A1 => n18471, A2 => n16645, B1 => n16881, B2 => 
                           n16648, ZN => n3928);
   U15541 : NAND2_X1 port map( A1 => n16719, A2 => n16673, ZN => n16650);
   U15542 : CLKBUF_X2 port map( A => n16650, Z => n16652);
   U15543 : NAND2_X1 port map( A1 => n13731, A2 => n16652, ZN => n16651);
   U15544 : OAI22_X1 port map( A1 => n16887, A2 => n16651, B1 => n16745, B2 => 
                           n16652, ZN => n3927);
   U15545 : CLKBUF_X2 port map( A => n16651, Z => n16649);
   U15546 : OAI22_X1 port map( A1 => n18120, A2 => n16649, B1 => n16816, B2 => 
                           n16650, ZN => n3926);
   U15547 : OAI22_X1 port map( A1 => n18804, A2 => n16651, B1 => n16817, B2 => 
                           n16652, ZN => n3925);
   U15548 : OAI22_X1 port map( A1 => n18805, A2 => n16649, B1 => n16818, B2 => 
                           n16650, ZN => n3924);
   U15549 : OAI22_X1 port map( A1 => n18121, A2 => n16649, B1 => n16819, B2 => 
                           n16650, ZN => n3923);
   U15550 : OAI22_X1 port map( A1 => n18122, A2 => n16649, B1 => n16820, B2 => 
                           n16652, ZN => n3922);
   U15551 : OAI22_X1 port map( A1 => n18472, A2 => n16649, B1 => n16821, B2 => 
                           n16650, ZN => n3921);
   U15552 : OAI22_X1 port map( A1 => n18123, A2 => n16649, B1 => n16822, B2 => 
                           n16652, ZN => n3920);
   U15553 : OAI22_X1 port map( A1 => n18473, A2 => n16649, B1 => n16823, B2 => 
                           n16652, ZN => n3919);
   U15554 : OAI22_X1 port map( A1 => n18474, A2 => n16649, B1 => n16824, B2 => 
                           n16652, ZN => n3918);
   U15555 : OAI22_X1 port map( A1 => n18475, A2 => n16649, B1 => n16825, B2 => 
                           n16652, ZN => n3917);
   U15556 : OAI22_X1 port map( A1 => n18806, A2 => n16649, B1 => n16826, B2 => 
                           n16652, ZN => n3916);
   U15557 : OAI22_X1 port map( A1 => n18124, A2 => n16651, B1 => n16827, B2 => 
                           n16650, ZN => n3915);
   U15558 : OAI22_X1 port map( A1 => n18125, A2 => n16649, B1 => n16828, B2 => 
                           n16650, ZN => n3914);
   U15559 : OAI22_X1 port map( A1 => n18476, A2 => n16649, B1 => n16829, B2 => 
                           n16650, ZN => n3913);
   U15560 : OAI22_X1 port map( A1 => n18126, A2 => n16651, B1 => n16830, B2 => 
                           n16652, ZN => n3912);
   U15561 : OAI22_X1 port map( A1 => n18127, A2 => n16651, B1 => n16831, B2 => 
                           n16650, ZN => n3911);
   U15562 : OAI22_X1 port map( A1 => n18477, A2 => n16649, B1 => n16832, B2 => 
                           n16650, ZN => n3910);
   U15563 : OAI22_X1 port map( A1 => n18478, A2 => n16649, B1 => n16833, B2 => 
                           n16650, ZN => n3909);
   U15564 : OAI22_X1 port map( A1 => n18479, A2 => n16651, B1 => n16834, B2 => 
                           n16652, ZN => n3908);
   U15565 : OAI22_X1 port map( A1 => n18480, A2 => n16651, B1 => n16835, B2 => 
                           n16650, ZN => n3907);
   U15566 : OAI22_X1 port map( A1 => n18128, A2 => n16649, B1 => n16836, B2 => 
                           n16652, ZN => n3906);
   U15567 : OAI22_X1 port map( A1 => n18481, A2 => n16649, B1 => n16837, B2 => 
                           n16652, ZN => n3905);
   U15568 : OAI22_X1 port map( A1 => n18482, A2 => n16649, B1 => n16838, B2 => 
                           n16650, ZN => n3904);
   U15569 : OAI22_X1 port map( A1 => n18483, A2 => n16649, B1 => n16839, B2 => 
                           n16652, ZN => n3903);
   U15570 : OAI22_X1 port map( A1 => n18129, A2 => n16651, B1 => n16840, B2 => 
                           n16650, ZN => n3902);
   U15571 : OAI22_X1 port map( A1 => n18484, A2 => n16649, B1 => n16841, B2 => 
                           n16650, ZN => n3901);
   U15572 : OAI22_X1 port map( A1 => n18485, A2 => n16651, B1 => n16842, B2 => 
                           n16650, ZN => n3900);
   U15573 : OAI22_X1 port map( A1 => n18130, A2 => n16649, B1 => n16843, B2 => 
                           n16650, ZN => n3899);
   U15574 : OAI22_X1 port map( A1 => n18486, A2 => n16651, B1 => n16844, B2 => 
                           n16650, ZN => n3898);
   U15575 : OAI22_X1 port map( A1 => n18487, A2 => n16649, B1 => n16845, B2 => 
                           n16650, ZN => n3897);
   U15576 : OAI22_X1 port map( A1 => n18488, A2 => n16651, B1 => n16846, B2 => 
                           n16650, ZN => n3896);
   U15577 : OAI22_X1 port map( A1 => n18489, A2 => n16649, B1 => n16847, B2 => 
                           n16650, ZN => n3895);
   U15578 : OAI22_X1 port map( A1 => n18131, A2 => n16651, B1 => n16848, B2 => 
                           n16650, ZN => n3894);
   U15579 : OAI22_X1 port map( A1 => n18132, A2 => n16649, B1 => n16849, B2 => 
                           n16650, ZN => n3893);
   U15580 : OAI22_X1 port map( A1 => n18490, A2 => n16651, B1 => n16850, B2 => 
                           n16652, ZN => n3892);
   U15581 : OAI22_X1 port map( A1 => n17823, A2 => n16651, B1 => n16851, B2 => 
                           n16652, ZN => n3891);
   U15582 : OAI22_X1 port map( A1 => n17451, A2 => n16649, B1 => n16852, B2 => 
                           n16652, ZN => n3890);
   U15583 : OAI22_X1 port map( A1 => n17212, A2 => n16651, B1 => n16853, B2 => 
                           n16652, ZN => n3889);
   U15584 : OAI22_X1 port map( A1 => n17213, A2 => n16649, B1 => n16854, B2 => 
                           n16652, ZN => n3888);
   U15585 : OAI22_X1 port map( A1 => n17452, A2 => n16651, B1 => n16855, B2 => 
                           n16652, ZN => n3887);
   U15586 : OAI22_X1 port map( A1 => n17214, A2 => n16649, B1 => n16856, B2 => 
                           n16652, ZN => n3886);
   U15587 : OAI22_X1 port map( A1 => n17453, A2 => n16649, B1 => n16857, B2 => 
                           n16652, ZN => n3885);
   U15588 : OAI22_X1 port map( A1 => n17215, A2 => n16649, B1 => n16858, B2 => 
                           n16652, ZN => n3884);
   U15589 : OAI22_X1 port map( A1 => n17454, A2 => n16649, B1 => n16859, B2 => 
                           n16652, ZN => n3883);
   U15590 : OAI22_X1 port map( A1 => n17216, A2 => n16649, B1 => n16860, B2 => 
                           n16652, ZN => n3882);
   U15591 : OAI22_X1 port map( A1 => n17217, A2 => n16649, B1 => n16861, B2 => 
                           n16652, ZN => n3881);
   U15592 : OAI22_X1 port map( A1 => n17218, A2 => n16649, B1 => n16862, B2 => 
                           n16652, ZN => n3880);
   U15593 : OAI22_X1 port map( A1 => n18491, A2 => n16651, B1 => n16863, B2 => 
                           n16652, ZN => n3879);
   U15594 : OAI22_X1 port map( A1 => n18492, A2 => n16651, B1 => n16864, B2 => 
                           n16652, ZN => n3878);
   U15595 : OAI22_X1 port map( A1 => n18133, A2 => n16649, B1 => n16865, B2 => 
                           n16652, ZN => n3877);
   U15596 : OAI22_X1 port map( A1 => n18493, A2 => n16649, B1 => n16866, B2 => 
                           n16652, ZN => n3876);
   U15597 : OAI22_X1 port map( A1 => n18134, A2 => n16651, B1 => n16867, B2 => 
                           n16652, ZN => n3875);
   U15598 : OAI22_X1 port map( A1 => n18135, A2 => n16649, B1 => n16868, B2 => 
                           n16652, ZN => n3874);
   U15599 : OAI22_X1 port map( A1 => n18136, A2 => n16651, B1 => n16869, B2 => 
                           n16652, ZN => n3873);
   U15600 : OAI22_X1 port map( A1 => n18494, A2 => n16649, B1 => n16870, B2 => 
                           n16652, ZN => n3872);
   U15601 : OAI22_X1 port map( A1 => n18137, A2 => n16651, B1 => n16871, B2 => 
                           n16652, ZN => n3871);
   U15602 : OAI22_X1 port map( A1 => n18138, A2 => n16651, B1 => n16872, B2 => 
                           n16652, ZN => n3870);
   U15603 : OAI22_X1 port map( A1 => n18495, A2 => n16649, B1 => n16873, B2 => 
                           n16652, ZN => n3869);
   U15604 : OAI22_X1 port map( A1 => n18807, A2 => n16649, B1 => n16874, B2 => 
                           n16650, ZN => n3868);
   U15605 : OAI22_X1 port map( A1 => n18139, A2 => n16651, B1 => n16875, B2 => 
                           n16652, ZN => n3867);
   U15606 : OAI22_X1 port map( A1 => n18140, A2 => n16649, B1 => n16876, B2 => 
                           n16652, ZN => n3866);
   U15607 : OAI22_X1 port map( A1 => n18141, A2 => n16651, B1 => n16878, B2 => 
                           n16650, ZN => n3865);
   U15608 : OAI22_X1 port map( A1 => n18142, A2 => n16649, B1 => n16881, B2 => 
                           n16652, ZN => n3864);
   U15609 : NAND2_X1 port map( A1 => n16724, A2 => n16673, ZN => n16654);
   U15610 : CLKBUF_X2 port map( A => n16654, Z => n16656);
   U15611 : NAND2_X1 port map( A1 => n13731, A2 => n16656, ZN => n16655);
   U15612 : OAI22_X1 port map( A1 => n16888, A2 => n16655, B1 => n16815, B2 => 
                           n16656, ZN => n3863);
   U15613 : CLKBUF_X2 port map( A => n16655, Z => n16653);
   U15614 : OAI22_X1 port map( A1 => n18496, A2 => n16653, B1 => n16746, B2 => 
                           n16654, ZN => n3862);
   U15615 : OAI22_X1 port map( A1 => n18143, A2 => n16655, B1 => n16747, B2 => 
                           n16656, ZN => n3861);
   U15616 : OAI22_X1 port map( A1 => n18144, A2 => n16653, B1 => n16748, B2 => 
                           n16654, ZN => n3860);
   U15617 : OAI22_X1 port map( A1 => n18145, A2 => n16653, B1 => n16749, B2 => 
                           n16654, ZN => n3859);
   U15618 : OAI22_X1 port map( A1 => n18146, A2 => n16653, B1 => n16750, B2 => 
                           n16656, ZN => n3858);
   U15619 : OAI22_X1 port map( A1 => n18147, A2 => n16653, B1 => n16751, B2 => 
                           n16654, ZN => n3857);
   U15620 : OAI22_X1 port map( A1 => n18148, A2 => n16653, B1 => n16752, B2 => 
                           n16656, ZN => n3856);
   U15621 : OAI22_X1 port map( A1 => n18497, A2 => n16653, B1 => n16753, B2 => 
                           n16656, ZN => n3855);
   U15622 : OAI22_X1 port map( A1 => n18498, A2 => n16653, B1 => n16754, B2 => 
                           n16656, ZN => n3854);
   U15623 : OAI22_X1 port map( A1 => n18149, A2 => n16653, B1 => n16755, B2 => 
                           n16656, ZN => n3853);
   U15624 : OAI22_X1 port map( A1 => n18499, A2 => n16653, B1 => n16756, B2 => 
                           n16656, ZN => n3852);
   U15625 : OAI22_X1 port map( A1 => n18150, A2 => n16655, B1 => n16757, B2 => 
                           n16654, ZN => n3851);
   U15626 : OAI22_X1 port map( A1 => n18500, A2 => n16653, B1 => n16758, B2 => 
                           n16654, ZN => n3850);
   U15627 : OAI22_X1 port map( A1 => n18151, A2 => n16653, B1 => n16759, B2 => 
                           n16654, ZN => n3849);
   U15628 : OAI22_X1 port map( A1 => n18501, A2 => n16655, B1 => n16760, B2 => 
                           n16656, ZN => n3848);
   U15629 : OAI22_X1 port map( A1 => n18502, A2 => n16655, B1 => n16761, B2 => 
                           n16654, ZN => n3847);
   U15630 : OAI22_X1 port map( A1 => n18503, A2 => n16653, B1 => n16762, B2 => 
                           n16654, ZN => n3846);
   U15631 : OAI22_X1 port map( A1 => n18504, A2 => n16653, B1 => n16763, B2 => 
                           n16654, ZN => n3845);
   U15632 : OAI22_X1 port map( A1 => n18808, A2 => n16655, B1 => n16764, B2 => 
                           n16656, ZN => n3844);
   U15633 : OAI22_X1 port map( A1 => n18505, A2 => n16655, B1 => n16765, B2 => 
                           n16654, ZN => n3843);
   U15634 : OAI22_X1 port map( A1 => n18506, A2 => n16653, B1 => n16766, B2 => 
                           n16656, ZN => n3842);
   U15635 : OAI22_X1 port map( A1 => n18809, A2 => n16653, B1 => n16767, B2 => 
                           n16656, ZN => n3841);
   U15636 : OAI22_X1 port map( A1 => n18152, A2 => n16653, B1 => n16768, B2 => 
                           n16654, ZN => n3840);
   U15637 : OAI22_X1 port map( A1 => n18507, A2 => n16653, B1 => n16769, B2 => 
                           n16656, ZN => n3839);
   U15638 : OAI22_X1 port map( A1 => n18508, A2 => n16655, B1 => n16770, B2 => 
                           n16654, ZN => n3838);
   U15639 : OAI22_X1 port map( A1 => n18509, A2 => n16653, B1 => n16771, B2 => 
                           n16654, ZN => n3837);
   U15640 : OAI22_X1 port map( A1 => n18510, A2 => n16655, B1 => n16772, B2 => 
                           n16654, ZN => n3836);
   U15641 : OAI22_X1 port map( A1 => n18153, A2 => n16653, B1 => n16773, B2 => 
                           n16654, ZN => n3835);
   U15642 : OAI22_X1 port map( A1 => n18511, A2 => n16655, B1 => n16774, B2 => 
                           n16654, ZN => n3834);
   U15643 : OAI22_X1 port map( A1 => n18512, A2 => n16653, B1 => n16775, B2 => 
                           n16654, ZN => n3833);
   U15644 : OAI22_X1 port map( A1 => n18810, A2 => n16655, B1 => n16776, B2 => 
                           n16654, ZN => n3832);
   U15645 : OAI22_X1 port map( A1 => n18154, A2 => n16653, B1 => n16777, B2 => 
                           n16654, ZN => n3831);
   U15646 : OAI22_X1 port map( A1 => n18513, A2 => n16655, B1 => n16778, B2 => 
                           n16654, ZN => n3830);
   U15647 : OAI22_X1 port map( A1 => n18155, A2 => n16653, B1 => n16779, B2 => 
                           n16654, ZN => n3829);
   U15648 : OAI22_X1 port map( A1 => n18514, A2 => n16655, B1 => n16781, B2 => 
                           n16656, ZN => n3828);
   U15649 : OAI22_X1 port map( A1 => n17219, A2 => n16655, B1 => n16782, B2 => 
                           n16656, ZN => n3827);
   U15650 : OAI22_X1 port map( A1 => n17220, A2 => n16653, B1 => n16783, B2 => 
                           n16656, ZN => n3826);
   U15651 : OAI22_X1 port map( A1 => n17824, A2 => n16655, B1 => n16784, B2 => 
                           n16656, ZN => n3825);
   U15652 : OAI22_X1 port map( A1 => n17221, A2 => n16653, B1 => n16785, B2 => 
                           n16656, ZN => n3824);
   U15653 : OAI22_X1 port map( A1 => n17455, A2 => n16655, B1 => n16786, B2 => 
                           n16656, ZN => n3823);
   U15654 : OAI22_X1 port map( A1 => n17825, A2 => n16653, B1 => n16787, B2 => 
                           n16656, ZN => n3822);
   U15655 : OAI22_X1 port map( A1 => n17826, A2 => n16653, B1 => n16788, B2 => 
                           n16656, ZN => n3821);
   U15656 : OAI22_X1 port map( A1 => n17456, A2 => n16653, B1 => n16789, B2 => 
                           n16656, ZN => n3820);
   U15657 : OAI22_X1 port map( A1 => n17457, A2 => n16653, B1 => n16790, B2 => 
                           n16656, ZN => n3819);
   U15658 : OAI22_X1 port map( A1 => n17458, A2 => n16653, B1 => n16791, B2 => 
                           n16656, ZN => n3818);
   U15659 : OAI22_X1 port map( A1 => n17459, A2 => n16653, B1 => n16792, B2 => 
                           n16656, ZN => n3817);
   U15660 : OAI22_X1 port map( A1 => n17222, A2 => n16653, B1 => n16793, B2 => 
                           n16656, ZN => n3816);
   U15661 : OAI22_X1 port map( A1 => n18156, A2 => n16655, B1 => n16794, B2 => 
                           n16656, ZN => n3815);
   U15662 : OAI22_X1 port map( A1 => n18515, A2 => n16655, B1 => n16795, B2 => 
                           n16656, ZN => n3814);
   U15663 : OAI22_X1 port map( A1 => n18516, A2 => n16653, B1 => n16796, B2 => 
                           n16656, ZN => n3813);
   U15664 : OAI22_X1 port map( A1 => n18517, A2 => n16653, B1 => n16797, B2 => 
                           n16656, ZN => n3812);
   U15665 : OAI22_X1 port map( A1 => n18811, A2 => n16655, B1 => n16798, B2 => 
                           n16656, ZN => n3811);
   U15666 : OAI22_X1 port map( A1 => n18157, A2 => n16653, B1 => n16799, B2 => 
                           n16656, ZN => n3810);
   U15667 : OAI22_X1 port map( A1 => n18158, A2 => n16655, B1 => n16800, B2 => 
                           n16656, ZN => n3809);
   U15668 : OAI22_X1 port map( A1 => n18518, A2 => n16653, B1 => n16801, B2 => 
                           n16656, ZN => n3808);
   U15669 : OAI22_X1 port map( A1 => n18519, A2 => n16655, B1 => n16802, B2 => 
                           n16656, ZN => n3807);
   U15670 : OAI22_X1 port map( A1 => n18520, A2 => n16655, B1 => n16803, B2 => 
                           n16656, ZN => n3806);
   U15671 : OAI22_X1 port map( A1 => n18812, A2 => n16653, B1 => n16804, B2 => 
                           n16656, ZN => n3805);
   U15672 : OAI22_X1 port map( A1 => n18159, A2 => n16653, B1 => n16805, B2 => 
                           n16654, ZN => n3804);
   U15673 : OAI22_X1 port map( A1 => n18160, A2 => n16655, B1 => n16806, B2 => 
                           n16656, ZN => n3803);
   U15674 : OAI22_X1 port map( A1 => n18521, A2 => n16653, B1 => n16808, B2 => 
                           n16656, ZN => n3802);
   U15675 : OAI22_X1 port map( A1 => n18161, A2 => n16655, B1 => n16810, B2 => 
                           n16654, ZN => n3801);
   U15676 : OAI22_X1 port map( A1 => n18522, A2 => n16653, B1 => n16812, B2 => 
                           n16656, ZN => n3800);
   U15677 : NAND2_X1 port map( A1 => n16729, A2 => n16673, ZN => n16657);
   U15678 : CLKBUF_X2 port map( A => n16657, Z => n16659);
   U15679 : NAND2_X1 port map( A1 => n13731, A2 => n16659, ZN => n16658);
   U15680 : OAI22_X1 port map( A1 => n16965, A2 => n16658, B1 => n16815, B2 => 
                           n16659, ZN => n3799);
   U15681 : OAI22_X1 port map( A1 => n18523, A2 => n16660, B1 => n16816, B2 => 
                           n16657, ZN => n3798);
   U15682 : OAI22_X1 port map( A1 => n18813, A2 => n16658, B1 => n16817, B2 => 
                           n16659, ZN => n3797);
   U15683 : OAI22_X1 port map( A1 => n18162, A2 => n16660, B1 => n16818, B2 => 
                           n16657, ZN => n3796);
   U15684 : OAI22_X1 port map( A1 => n18814, A2 => n16660, B1 => n16819, B2 => 
                           n16657, ZN => n3795);
   U15685 : OAI22_X1 port map( A1 => n18163, A2 => n16658, B1 => n16820, B2 => 
                           n16659, ZN => n3794);
   U15686 : OAI22_X1 port map( A1 => n18524, A2 => n16660, B1 => n16821, B2 => 
                           n16657, ZN => n3793);
   U15687 : OAI22_X1 port map( A1 => n18815, A2 => n16658, B1 => n16822, B2 => 
                           n16659, ZN => n3792);
   U15688 : OAI22_X1 port map( A1 => n18816, A2 => n16660, B1 => n16823, B2 => 
                           n16659, ZN => n3791);
   U15689 : OAI22_X1 port map( A1 => n18164, A2 => n16658, B1 => n16824, B2 => 
                           n16659, ZN => n3790);
   U15690 : OAI22_X1 port map( A1 => n18525, A2 => n16660, B1 => n16825, B2 => 
                           n16659, ZN => n3789);
   U15691 : OAI22_X1 port map( A1 => n18165, A2 => n16660, B1 => n16826, B2 => 
                           n16659, ZN => n3788);
   U15692 : OAI22_X1 port map( A1 => n18526, A2 => n16658, B1 => n16827, B2 => 
                           n16657, ZN => n3787);
   U15693 : OAI22_X1 port map( A1 => n18527, A2 => n16660, B1 => n16828, B2 => 
                           n16657, ZN => n3786);
   U15694 : OAI22_X1 port map( A1 => n18166, A2 => n16660, B1 => n16829, B2 => 
                           n16657, ZN => n3785);
   U15695 : OAI22_X1 port map( A1 => n18528, A2 => n16658, B1 => n16830, B2 => 
                           n16659, ZN => n3784);
   U15696 : OAI22_X1 port map( A1 => n18529, A2 => n16658, B1 => n16831, B2 => 
                           n16657, ZN => n3783);
   U15697 : OAI22_X1 port map( A1 => n18530, A2 => n16660, B1 => n16832, B2 => 
                           n16657, ZN => n3782);
   U15698 : OAI22_X1 port map( A1 => n18531, A2 => n16660, B1 => n16833, B2 => 
                           n16657, ZN => n3781);
   U15699 : OAI22_X1 port map( A1 => n18167, A2 => n16658, B1 => n16834, B2 => 
                           n16659, ZN => n3780);
   U15700 : OAI22_X1 port map( A1 => n18817, A2 => n16658, B1 => n16835, B2 => 
                           n16657, ZN => n3779);
   U15701 : OAI22_X1 port map( A1 => n18532, A2 => n16660, B1 => n16836, B2 => 
                           n16659, ZN => n3778);
   U15702 : OAI22_X1 port map( A1 => n18818, A2 => n16660, B1 => n16837, B2 => 
                           n16659, ZN => n3777);
   U15703 : OAI22_X1 port map( A1 => n18168, A2 => n16660, B1 => n16838, B2 => 
                           n16657, ZN => n3776);
   U15704 : OAI22_X1 port map( A1 => n18533, A2 => n16660, B1 => n16839, B2 => 
                           n16659, ZN => n3775);
   U15705 : OAI22_X1 port map( A1 => n18819, A2 => n16658, B1 => n16840, B2 => 
                           n16657, ZN => n3774);
   U15706 : OAI22_X1 port map( A1 => n18534, A2 => n16660, B1 => n16841, B2 => 
                           n16657, ZN => n3773);
   U15707 : OAI22_X1 port map( A1 => n18169, A2 => n16658, B1 => n16842, B2 => 
                           n16657, ZN => n3772);
   U15708 : OAI22_X1 port map( A1 => n18535, A2 => n16660, B1 => n16843, B2 => 
                           n16657, ZN => n3771);
   U15709 : OAI22_X1 port map( A1 => n18536, A2 => n16658, B1 => n16844, B2 => 
                           n16657, ZN => n3770);
   U15710 : OAI22_X1 port map( A1 => n18820, A2 => n16660, B1 => n16845, B2 => 
                           n16657, ZN => n3769);
   U15711 : OAI22_X1 port map( A1 => n18170, A2 => n16658, B1 => n16846, B2 => 
                           n16657, ZN => n3768);
   U15712 : OAI22_X1 port map( A1 => n18821, A2 => n16660, B1 => n16847, B2 => 
                           n16657, ZN => n3767);
   U15713 : OAI22_X1 port map( A1 => n18171, A2 => n16658, B1 => n16848, B2 => 
                           n16657, ZN => n3766);
   U15714 : OAI22_X1 port map( A1 => n18822, A2 => n16660, B1 => n16849, B2 => 
                           n16657, ZN => n3765);
   U15715 : OAI22_X1 port map( A1 => n18172, A2 => n16658, B1 => n16850, B2 => 
                           n16659, ZN => n3764);
   U15716 : CLKBUF_X2 port map( A => n16658, Z => n16660);
   U15717 : OAI22_X1 port map( A1 => n17223, A2 => n16660, B1 => n16851, B2 => 
                           n16659, ZN => n3763);
   U15718 : OAI22_X1 port map( A1 => n17460, A2 => n16660, B1 => n16852, B2 => 
                           n16659, ZN => n3762);
   U15719 : OAI22_X1 port map( A1 => n17461, A2 => n16660, B1 => n16853, B2 => 
                           n16659, ZN => n3761);
   U15720 : OAI22_X1 port map( A1 => n17827, A2 => n16660, B1 => n16854, B2 => 
                           n16659, ZN => n3760);
   U15721 : OAI22_X1 port map( A1 => n17828, A2 => n16660, B1 => n16855, B2 => 
                           n16659, ZN => n3759);
   U15722 : OAI22_X1 port map( A1 => n17462, A2 => n16660, B1 => n16856, B2 => 
                           n16659, ZN => n3758);
   U15723 : OAI22_X1 port map( A1 => n17829, A2 => n16660, B1 => n16857, B2 => 
                           n16659, ZN => n3757);
   U15724 : OAI22_X1 port map( A1 => n17224, A2 => n16660, B1 => n16858, B2 => 
                           n16659, ZN => n3756);
   U15725 : OAI22_X1 port map( A1 => n17463, A2 => n16660, B1 => n16859, B2 => 
                           n16659, ZN => n3755);
   U15726 : OAI22_X1 port map( A1 => n17464, A2 => n16660, B1 => n16860, B2 => 
                           n16659, ZN => n3754);
   U15727 : OAI22_X1 port map( A1 => n17225, A2 => n16660, B1 => n16861, B2 => 
                           n16659, ZN => n3753);
   U15728 : OAI22_X1 port map( A1 => n17465, A2 => n16660, B1 => n16862, B2 => 
                           n16659, ZN => n3752);
   U15729 : OAI22_X1 port map( A1 => n18173, A2 => n16658, B1 => n16863, B2 => 
                           n16659, ZN => n3751);
   U15730 : OAI22_X1 port map( A1 => n18174, A2 => n16658, B1 => n16864, B2 => 
                           n16659, ZN => n3750);
   U15731 : OAI22_X1 port map( A1 => n18537, A2 => n16660, B1 => n16865, B2 => 
                           n16659, ZN => n3749);
   U15732 : OAI22_X1 port map( A1 => n18823, A2 => n16660, B1 => n16866, B2 => 
                           n16659, ZN => n3748);
   U15733 : OAI22_X1 port map( A1 => n18538, A2 => n16658, B1 => n16867, B2 => 
                           n16659, ZN => n3747);
   U15734 : OAI22_X1 port map( A1 => n18824, A2 => n16660, B1 => n16868, B2 => 
                           n16659, ZN => n3746);
   U15735 : OAI22_X1 port map( A1 => n18825, A2 => n16658, B1 => n16869, B2 => 
                           n16659, ZN => n3745);
   U15736 : OAI22_X1 port map( A1 => n18826, A2 => n16660, B1 => n16870, B2 => 
                           n16659, ZN => n3744);
   U15737 : OAI22_X1 port map( A1 => n18827, A2 => n16658, B1 => n16871, B2 => 
                           n16659, ZN => n3743);
   U15738 : OAI22_X1 port map( A1 => n18175, A2 => n16658, B1 => n16872, B2 => 
                           n16659, ZN => n3742);
   U15739 : OAI22_X1 port map( A1 => n18828, A2 => n16660, B1 => n16873, B2 => 
                           n16659, ZN => n3741);
   U15740 : OAI22_X1 port map( A1 => n18539, A2 => n16660, B1 => n16874, B2 => 
                           n16657, ZN => n3740);
   U15741 : OAI22_X1 port map( A1 => n18540, A2 => n16658, B1 => n16875, B2 => 
                           n16659, ZN => n3739);
   U15742 : OAI22_X1 port map( A1 => n18541, A2 => n16660, B1 => n16876, B2 => 
                           n16659, ZN => n3738);
   U15743 : OAI22_X1 port map( A1 => n18829, A2 => n16658, B1 => n16878, B2 => 
                           n16657, ZN => n3737);
   U15744 : OAI22_X1 port map( A1 => n18176, A2 => n16660, B1 => n16881, B2 => 
                           n16659, ZN => n3736);
   U15745 : NAND2_X1 port map( A1 => n16734, A2 => n16673, ZN => n16663);
   U15746 : NAND2_X1 port map( A1 => n13731, A2 => n16662, ZN => n16664);
   U15747 : OAI22_X1 port map( A1 => n17226, A2 => n16664, B1 => n16745, B2 => 
                           n16663, ZN => n3735);
   U15748 : CLKBUF_X2 port map( A => n16664, Z => n16661);
   U15749 : CLKBUF_X2 port map( A => n16663, Z => n16662);
   U15750 : OAI22_X1 port map( A1 => n17227, A2 => n16661, B1 => n16746, B2 => 
                           n16662, ZN => n3734);
   U15751 : OAI22_X1 port map( A1 => n17228, A2 => n16664, B1 => n16747, B2 => 
                           n16663, ZN => n3733);
   U15752 : OAI22_X1 port map( A1 => n17466, A2 => n16661, B1 => n16748, B2 => 
                           n16663, ZN => n3732);
   U15753 : OAI22_X1 port map( A1 => n17467, A2 => n16661, B1 => n16749, B2 => 
                           n16663, ZN => n3731);
   U15754 : OAI22_X1 port map( A1 => n17468, A2 => n16661, B1 => n16750, B2 => 
                           n16663, ZN => n3730);
   U15755 : OAI22_X1 port map( A1 => n17469, A2 => n16661, B1 => n16751, B2 => 
                           n16662, ZN => n3729);
   U15756 : OAI22_X1 port map( A1 => n17470, A2 => n16661, B1 => n16752, B2 => 
                           n16663, ZN => n3728);
   U15757 : OAI22_X1 port map( A1 => n17471, A2 => n16661, B1 => n16753, B2 => 
                           n16662, ZN => n3727);
   U15758 : OAI22_X1 port map( A1 => n17830, A2 => n16661, B1 => n16754, B2 => 
                           n16663, ZN => n3726);
   U15759 : OAI22_X1 port map( A1 => n17472, A2 => n16661, B1 => n16755, B2 => 
                           n16662, ZN => n3725);
   U15760 : OAI22_X1 port map( A1 => n17473, A2 => n16661, B1 => n16756, B2 => 
                           n16662, ZN => n3724);
   U15761 : OAI22_X1 port map( A1 => n18542, A2 => n16664, B1 => n16757, B2 => 
                           n16663, ZN => n3723);
   U15762 : OAI22_X1 port map( A1 => n18543, A2 => n16661, B1 => n16758, B2 => 
                           n16662, ZN => n3722);
   U15763 : OAI22_X1 port map( A1 => n18177, A2 => n16661, B1 => n16759, B2 => 
                           n16663, ZN => n3721);
   U15764 : OAI22_X1 port map( A1 => n18830, A2 => n16664, B1 => n16760, B2 => 
                           n16662, ZN => n3720);
   U15765 : OAI22_X1 port map( A1 => n18178, A2 => n16664, B1 => n16761, B2 => 
                           n16663, ZN => n3719);
   U15766 : OAI22_X1 port map( A1 => n18544, A2 => n16661, B1 => n16762, B2 => 
                           n16662, ZN => n3718);
   U15767 : OAI22_X1 port map( A1 => n18831, A2 => n16661, B1 => n16763, B2 => 
                           n16663, ZN => n3717);
   U15768 : OAI22_X1 port map( A1 => n18545, A2 => n16664, B1 => n16764, B2 => 
                           n16662, ZN => n3716);
   U15769 : OAI22_X1 port map( A1 => n18546, A2 => n16664, B1 => n16765, B2 => 
                           n16662, ZN => n3715);
   U15770 : OAI22_X1 port map( A1 => n18179, A2 => n16661, B1 => n16766, B2 => 
                           n16662, ZN => n3714);
   U15771 : OAI22_X1 port map( A1 => n18547, A2 => n16661, B1 => n16767, B2 => 
                           n16662, ZN => n3713);
   U15772 : OAI22_X1 port map( A1 => n18548, A2 => n16661, B1 => n16768, B2 => 
                           n16663, ZN => n3712);
   U15773 : OAI22_X1 port map( A1 => n18549, A2 => n16661, B1 => n16769, B2 => 
                           n16662, ZN => n3711);
   U15774 : OAI22_X1 port map( A1 => n18180, A2 => n16664, B1 => n16770, B2 => 
                           n16663, ZN => n3710);
   U15775 : OAI22_X1 port map( A1 => n18550, A2 => n16661, B1 => n16771, B2 => 
                           n16663, ZN => n3709);
   U15776 : OAI22_X1 port map( A1 => n18551, A2 => n16664, B1 => n16772, B2 => 
                           n16663, ZN => n3708);
   U15777 : OAI22_X1 port map( A1 => n18552, A2 => n16661, B1 => n16773, B2 => 
                           n16663, ZN => n3707);
   U15778 : OAI22_X1 port map( A1 => n18832, A2 => n16664, B1 => n16774, B2 => 
                           n16663, ZN => n3706);
   U15779 : OAI22_X1 port map( A1 => n18833, A2 => n16661, B1 => n16775, B2 => 
                           n16663, ZN => n3705);
   U15780 : OAI22_X1 port map( A1 => n18553, A2 => n16664, B1 => n16776, B2 => 
                           n16663, ZN => n3704);
   U15781 : OAI22_X1 port map( A1 => n18554, A2 => n16661, B1 => n16777, B2 => 
                           n16663, ZN => n3703);
   U15782 : OAI22_X1 port map( A1 => n18555, A2 => n16664, B1 => n16778, B2 => 
                           n16663, ZN => n3702);
   U15783 : OAI22_X1 port map( A1 => n18834, A2 => n16661, B1 => n16779, B2 => 
                           n16663, ZN => n3701);
   U15784 : OAI22_X1 port map( A1 => n18556, A2 => n16664, B1 => n16781, B2 => 
                           n16662, ZN => n3700);
   U15785 : OAI22_X1 port map( A1 => n17831, A2 => n16664, B1 => n16782, B2 => 
                           n16662, ZN => n3699);
   U15786 : OAI22_X1 port map( A1 => n17474, A2 => n16661, B1 => n16783, B2 => 
                           n16662, ZN => n3698);
   U15787 : OAI22_X1 port map( A1 => n17475, A2 => n16664, B1 => n16784, B2 => 
                           n16662, ZN => n3697);
   U15788 : OAI22_X1 port map( A1 => n17229, A2 => n16661, B1 => n16785, B2 => 
                           n16662, ZN => n3696);
   U15789 : OAI22_X1 port map( A1 => n17832, A2 => n16664, B1 => n16786, B2 => 
                           n16662, ZN => n3695);
   U15790 : OAI22_X1 port map( A1 => n17476, A2 => n16661, B1 => n16787, B2 => 
                           n16662, ZN => n3694);
   U15791 : OAI22_X1 port map( A1 => n17477, A2 => n16661, B1 => n16788, B2 => 
                           n16662, ZN => n3693);
   U15792 : OAI22_X1 port map( A1 => n17478, A2 => n16661, B1 => n16789, B2 => 
                           n16662, ZN => n3692);
   U15793 : OAI22_X1 port map( A1 => n17230, A2 => n16661, B1 => n16790, B2 => 
                           n16662, ZN => n3691);
   U15794 : OAI22_X1 port map( A1 => n17479, A2 => n16661, B1 => n16791, B2 => 
                           n16662, ZN => n3690);
   U15795 : OAI22_X1 port map( A1 => n17833, A2 => n16661, B1 => n16792, B2 => 
                           n16662, ZN => n3689);
   U15796 : OAI22_X1 port map( A1 => n17834, A2 => n16661, B1 => n16793, B2 => 
                           n16662, ZN => n3688);
   U15797 : OAI22_X1 port map( A1 => n18557, A2 => n16664, B1 => n16794, B2 => 
                           n16662, ZN => n3687);
   U15798 : OAI22_X1 port map( A1 => n18835, A2 => n16664, B1 => n16795, B2 => 
                           n16662, ZN => n3686);
   U15799 : OAI22_X1 port map( A1 => n18558, A2 => n16661, B1 => n16796, B2 => 
                           n16662, ZN => n3685);
   U15800 : OAI22_X1 port map( A1 => n18836, A2 => n16661, B1 => n16797, B2 => 
                           n16662, ZN => n3684);
   U15801 : OAI22_X1 port map( A1 => n18559, A2 => n16664, B1 => n16798, B2 => 
                           n16662, ZN => n3683);
   U15802 : OAI22_X1 port map( A1 => n18837, A2 => n16661, B1 => n16799, B2 => 
                           n16662, ZN => n3682);
   U15803 : OAI22_X1 port map( A1 => n18560, A2 => n16664, B1 => n16800, B2 => 
                           n16662, ZN => n3681);
   U15804 : OAI22_X1 port map( A1 => n18561, A2 => n16661, B1 => n16801, B2 => 
                           n16662, ZN => n3680);
   U15805 : OAI22_X1 port map( A1 => n18562, A2 => n16664, B1 => n16802, B2 => 
                           n16662, ZN => n3679);
   U15806 : OAI22_X1 port map( A1 => n18838, A2 => n16664, B1 => n16803, B2 => 
                           n16662, ZN => n3678);
   U15807 : OAI22_X1 port map( A1 => n18181, A2 => n16661, B1 => n16804, B2 => 
                           n16662, ZN => n3677);
   U15808 : OAI22_X1 port map( A1 => n18182, A2 => n16661, B1 => n16805, B2 => 
                           n16663, ZN => n3676);
   U15809 : OAI22_X1 port map( A1 => n18183, A2 => n16664, B1 => n16806, B2 => 
                           n16662, ZN => n3675);
   U15810 : OAI22_X1 port map( A1 => n18563, A2 => n16661, B1 => n16808, B2 => 
                           n16662, ZN => n3674);
   U15811 : OAI22_X1 port map( A1 => n18184, A2 => n16664, B1 => n16810, B2 => 
                           n16663, ZN => n3673);
   U15812 : OAI22_X1 port map( A1 => n18185, A2 => n16661, B1 => n16812, B2 => 
                           n16662, ZN => n3672);
   U15813 : NAND2_X1 port map( A1 => n16739, A2 => n16673, ZN => n16667);
   U15814 : NAND2_X1 port map( A1 => n13731, A2 => n16666, ZN => n16668);
   U15815 : OAI22_X1 port map( A1 => n17231, A2 => n16668, B1 => n16745, B2 => 
                           n16667, ZN => n3671);
   U15816 : CLKBUF_X2 port map( A => n16668, Z => n16665);
   U15817 : CLKBUF_X2 port map( A => n16667, Z => n16666);
   U15818 : OAI22_X1 port map( A1 => n17835, A2 => n16665, B1 => n16746, B2 => 
                           n16666, ZN => n3670);
   U15819 : OAI22_X1 port map( A1 => n17836, A2 => n16668, B1 => n16747, B2 => 
                           n16667, ZN => n3669);
   U15820 : OAI22_X1 port map( A1 => n17837, A2 => n16665, B1 => n16748, B2 => 
                           n16667, ZN => n3668);
   U15821 : OAI22_X1 port map( A1 => n17838, A2 => n16665, B1 => n16749, B2 => 
                           n16667, ZN => n3667);
   U15822 : OAI22_X1 port map( A1 => n17839, A2 => n16665, B1 => n16750, B2 => 
                           n16667, ZN => n3666);
   U15823 : OAI22_X1 port map( A1 => n17480, A2 => n16665, B1 => n16751, B2 => 
                           n16666, ZN => n3665);
   U15824 : OAI22_X1 port map( A1 => n17840, A2 => n16665, B1 => n16752, B2 => 
                           n16667, ZN => n3664);
   U15825 : OAI22_X1 port map( A1 => n17481, A2 => n16665, B1 => n16753, B2 => 
                           n16666, ZN => n3663);
   U15826 : OAI22_X1 port map( A1 => n17482, A2 => n16665, B1 => n16754, B2 => 
                           n16667, ZN => n3662);
   U15827 : OAI22_X1 port map( A1 => n17841, A2 => n16665, B1 => n16755, B2 => 
                           n16666, ZN => n3661);
   U15828 : OAI22_X1 port map( A1 => n17842, A2 => n16665, B1 => n16756, B2 => 
                           n16666, ZN => n3660);
   U15829 : OAI22_X1 port map( A1 => n18564, A2 => n16668, B1 => n16757, B2 => 
                           n16667, ZN => n3659);
   U15830 : OAI22_X1 port map( A1 => n18839, A2 => n16665, B1 => n16758, B2 => 
                           n16666, ZN => n3658);
   U15831 : OAI22_X1 port map( A1 => n18840, A2 => n16665, B1 => n16759, B2 => 
                           n16667, ZN => n3657);
   U15832 : OAI22_X1 port map( A1 => n18841, A2 => n16668, B1 => n16760, B2 => 
                           n16666, ZN => n3656);
   U15833 : OAI22_X1 port map( A1 => n18842, A2 => n16668, B1 => n16761, B2 => 
                           n16667, ZN => n3655);
   U15834 : OAI22_X1 port map( A1 => n18843, A2 => n16665, B1 => n16762, B2 => 
                           n16666, ZN => n3654);
   U15835 : OAI22_X1 port map( A1 => n18844, A2 => n16665, B1 => n16763, B2 => 
                           n16667, ZN => n3653);
   U15836 : OAI22_X1 port map( A1 => n18565, A2 => n16668, B1 => n16764, B2 => 
                           n16666, ZN => n3652);
   U15837 : OAI22_X1 port map( A1 => n18566, A2 => n16668, B1 => n16765, B2 => 
                           n16666, ZN => n3651);
   U15838 : OAI22_X1 port map( A1 => n18845, A2 => n16665, B1 => n16766, B2 => 
                           n16666, ZN => n3650);
   U15839 : OAI22_X1 port map( A1 => n18567, A2 => n16665, B1 => n16767, B2 => 
                           n16666, ZN => n3649);
   U15840 : OAI22_X1 port map( A1 => n18846, A2 => n16665, B1 => n16768, B2 => 
                           n16667, ZN => n3648);
   U15841 : OAI22_X1 port map( A1 => n18568, A2 => n16665, B1 => n16769, B2 => 
                           n16666, ZN => n3647);
   U15842 : OAI22_X1 port map( A1 => n18847, A2 => n16668, B1 => n16770, B2 => 
                           n16667, ZN => n3646);
   U15843 : OAI22_X1 port map( A1 => n18569, A2 => n16665, B1 => n16771, B2 => 
                           n16667, ZN => n3645);
   U15844 : OAI22_X1 port map( A1 => n18570, A2 => n16668, B1 => n16772, B2 => 
                           n16667, ZN => n3644);
   U15845 : OAI22_X1 port map( A1 => n18848, A2 => n16665, B1 => n16773, B2 => 
                           n16667, ZN => n3643);
   U15846 : OAI22_X1 port map( A1 => n18849, A2 => n16668, B1 => n16774, B2 => 
                           n16667, ZN => n3642);
   U15847 : OAI22_X1 port map( A1 => n18571, A2 => n16665, B1 => n16775, B2 => 
                           n16667, ZN => n3641);
   U15848 : OAI22_X1 port map( A1 => n18850, A2 => n16668, B1 => n16776, B2 => 
                           n16667, ZN => n3640);
   U15849 : OAI22_X1 port map( A1 => n18572, A2 => n16665, B1 => n16777, B2 => 
                           n16667, ZN => n3639);
   U15850 : OAI22_X1 port map( A1 => n18851, A2 => n16668, B1 => n16778, B2 => 
                           n16667, ZN => n3638);
   U15851 : OAI22_X1 port map( A1 => n18573, A2 => n16665, B1 => n16779, B2 => 
                           n16667, ZN => n3637);
   U15852 : OAI22_X1 port map( A1 => n18574, A2 => n16668, B1 => n16781, B2 => 
                           n16666, ZN => n3636);
   U15853 : OAI22_X1 port map( A1 => n17232, A2 => n16668, B1 => n16782, B2 => 
                           n16666, ZN => n3635);
   U15854 : OAI22_X1 port map( A1 => n17843, A2 => n16665, B1 => n16783, B2 => 
                           n16666, ZN => n3634);
   U15855 : OAI22_X1 port map( A1 => n17233, A2 => n16668, B1 => n16784, B2 => 
                           n16666, ZN => n3633);
   U15856 : OAI22_X1 port map( A1 => n17483, A2 => n16665, B1 => n16785, B2 => 
                           n16666, ZN => n3632);
   U15857 : OAI22_X1 port map( A1 => n17484, A2 => n16668, B1 => n16786, B2 => 
                           n16666, ZN => n3631);
   U15858 : OAI22_X1 port map( A1 => n17844, A2 => n16665, B1 => n16787, B2 => 
                           n16666, ZN => n3630);
   U15859 : OAI22_X1 port map( A1 => n17485, A2 => n16665, B1 => n16788, B2 => 
                           n16666, ZN => n3629);
   U15860 : OAI22_X1 port map( A1 => n17845, A2 => n16665, B1 => n16789, B2 => 
                           n16666, ZN => n3628);
   U15861 : OAI22_X1 port map( A1 => n17846, A2 => n16665, B1 => n16790, B2 => 
                           n16666, ZN => n3627);
   U15862 : OAI22_X1 port map( A1 => n17847, A2 => n16665, B1 => n16791, B2 => 
                           n16666, ZN => n3626);
   U15863 : OAI22_X1 port map( A1 => n17486, A2 => n16665, B1 => n16792, B2 => 
                           n16666, ZN => n3625);
   U15864 : OAI22_X1 port map( A1 => n17487, A2 => n16665, B1 => n16793, B2 => 
                           n16666, ZN => n3624);
   U15865 : OAI22_X1 port map( A1 => n18575, A2 => n16668, B1 => n16794, B2 => 
                           n16666, ZN => n3623);
   U15866 : OAI22_X1 port map( A1 => n18576, A2 => n16668, B1 => n16795, B2 => 
                           n16666, ZN => n3622);
   U15867 : OAI22_X1 port map( A1 => n18577, A2 => n16665, B1 => n16796, B2 => 
                           n16666, ZN => n3621);
   U15868 : OAI22_X1 port map( A1 => n18578, A2 => n16665, B1 => n16797, B2 => 
                           n16666, ZN => n3620);
   U15869 : OAI22_X1 port map( A1 => n18579, A2 => n16668, B1 => n16798, B2 => 
                           n16666, ZN => n3619);
   U15870 : OAI22_X1 port map( A1 => n18580, A2 => n16665, B1 => n16799, B2 => 
                           n16666, ZN => n3618);
   U15871 : OAI22_X1 port map( A1 => n18852, A2 => n16668, B1 => n16800, B2 => 
                           n16666, ZN => n3617);
   U15872 : OAI22_X1 port map( A1 => n18581, A2 => n16665, B1 => n16801, B2 => 
                           n16666, ZN => n3616);
   U15873 : OAI22_X1 port map( A1 => n18853, A2 => n16668, B1 => n16802, B2 => 
                           n16666, ZN => n3615);
   U15874 : OAI22_X1 port map( A1 => n18582, A2 => n16668, B1 => n16803, B2 => 
                           n16666, ZN => n3614);
   U15875 : OAI22_X1 port map( A1 => n18854, A2 => n16665, B1 => n16804, B2 => 
                           n16666, ZN => n3613);
   U15876 : OAI22_X1 port map( A1 => n18855, A2 => n16665, B1 => n16805, B2 => 
                           n16667, ZN => n3612);
   U15877 : OAI22_X1 port map( A1 => n18856, A2 => n16668, B1 => n16806, B2 => 
                           n16666, ZN => n3611);
   U15878 : OAI22_X1 port map( A1 => n18857, A2 => n16665, B1 => n16808, B2 => 
                           n16666, ZN => n3610);
   U15879 : OAI22_X1 port map( A1 => n18858, A2 => n16668, B1 => n16810, B2 => 
                           n16667, ZN => n3609);
   U15880 : OAI22_X1 port map( A1 => n18859, A2 => n16665, B1 => n16812, B2 => 
                           n16666, ZN => n3608);
   U15881 : NAND2_X1 port map( A1 => n16744, A2 => n16673, ZN => n16670);
   U15882 : CLKBUF_X2 port map( A => n16670, Z => n16672);
   U15883 : NAND2_X1 port map( A1 => n13731, A2 => n16672, ZN => n16671);
   U15884 : OAI22_X1 port map( A1 => n17171, A2 => n16671, B1 => n16745, B2 => 
                           n16670, ZN => n3607);
   U15885 : CLKBUF_X2 port map( A => n16671, Z => n16669);
   U15886 : OAI22_X1 port map( A1 => n17234, A2 => n16669, B1 => n16746, B2 => 
                           n16672, ZN => n3606);
   U15887 : OAI22_X1 port map( A1 => n17488, A2 => n16671, B1 => n16747, B2 => 
                           n16670, ZN => n3605);
   U15888 : OAI22_X1 port map( A1 => n17489, A2 => n16669, B1 => n16748, B2 => 
                           n16670, ZN => n3604);
   U15889 : OAI22_X1 port map( A1 => n17490, A2 => n16669, B1 => n16749, B2 => 
                           n16672, ZN => n3603);
   U15890 : OAI22_X1 port map( A1 => n17491, A2 => n16669, B1 => n16750, B2 => 
                           n16670, ZN => n3602);
   U15891 : OAI22_X1 port map( A1 => n17235, A2 => n16669, B1 => n16751, B2 => 
                           n16672, ZN => n3601);
   U15892 : OAI22_X1 port map( A1 => n17236, A2 => n16669, B1 => n16752, B2 => 
                           n16672, ZN => n3600);
   U15893 : OAI22_X1 port map( A1 => n17237, A2 => n16669, B1 => n16753, B2 => 
                           n16672, ZN => n3599);
   U15894 : OAI22_X1 port map( A1 => n17238, A2 => n16669, B1 => n16754, B2 => 
                           n16672, ZN => n3598);
   U15895 : OAI22_X1 port map( A1 => n17492, A2 => n16669, B1 => n16755, B2 => 
                           n16672, ZN => n3597);
   U15896 : OAI22_X1 port map( A1 => n17493, A2 => n16669, B1 => n16756, B2 => 
                           n16670, ZN => n3596);
   U15897 : OAI22_X1 port map( A1 => n18583, A2 => n16671, B1 => n16757, B2 => 
                           n16670, ZN => n3595);
   U15898 : OAI22_X1 port map( A1 => n18584, A2 => n16669, B1 => n16758, B2 => 
                           n16672, ZN => n3594);
   U15899 : OAI22_X1 port map( A1 => n18585, A2 => n16669, B1 => n16759, B2 => 
                           n16670, ZN => n3593);
   U15900 : OAI22_X1 port map( A1 => n18586, A2 => n16671, B1 => n16760, B2 => 
                           n16670, ZN => n3592);
   U15901 : OAI22_X1 port map( A1 => n18587, A2 => n16671, B1 => n16761, B2 => 
                           n16670, ZN => n3591);
   U15902 : OAI22_X1 port map( A1 => n18186, A2 => n16669, B1 => n16762, B2 => 
                           n16672, ZN => n3590);
   U15903 : OAI22_X1 port map( A1 => n18187, A2 => n16669, B1 => n16763, B2 => 
                           n16670, ZN => n3589);
   U15904 : OAI22_X1 port map( A1 => n18188, A2 => n16671, B1 => n16764, B2 => 
                           n16670, ZN => n3588);
   U15905 : OAI22_X1 port map( A1 => n18588, A2 => n16671, B1 => n16765, B2 => 
                           n16672, ZN => n3587);
   U15906 : OAI22_X1 port map( A1 => n18189, A2 => n16669, B1 => n16766, B2 => 
                           n16672, ZN => n3586);
   U15907 : OAI22_X1 port map( A1 => n18860, A2 => n16669, B1 => n16767, B2 => 
                           n16672, ZN => n3585);
   U15908 : OAI22_X1 port map( A1 => n18589, A2 => n16669, B1 => n16768, B2 => 
                           n16670, ZN => n3584);
   U15909 : OAI22_X1 port map( A1 => n18190, A2 => n16669, B1 => n16769, B2 => 
                           n16672, ZN => n3583);
   U15910 : OAI22_X1 port map( A1 => n18191, A2 => n16671, B1 => n16770, B2 => 
                           n16670, ZN => n3582);
   U15911 : OAI22_X1 port map( A1 => n18192, A2 => n16669, B1 => n16771, B2 => 
                           n16670, ZN => n3581);
   U15912 : OAI22_X1 port map( A1 => n18193, A2 => n16671, B1 => n16772, B2 => 
                           n16670, ZN => n3580);
   U15913 : OAI22_X1 port map( A1 => n18590, A2 => n16669, B1 => n16773, B2 => 
                           n16670, ZN => n3579);
   U15914 : OAI22_X1 port map( A1 => n18591, A2 => n16671, B1 => n16774, B2 => 
                           n16670, ZN => n3578);
   U15915 : OAI22_X1 port map( A1 => n18592, A2 => n16669, B1 => n16775, B2 => 
                           n16670, ZN => n3577);
   U15916 : OAI22_X1 port map( A1 => n18194, A2 => n16671, B1 => n16776, B2 => 
                           n16670, ZN => n3576);
   U15917 : OAI22_X1 port map( A1 => n18593, A2 => n16669, B1 => n16777, B2 => 
                           n16670, ZN => n3575);
   U15918 : OAI22_X1 port map( A1 => n18195, A2 => n16671, B1 => n16778, B2 => 
                           n16670, ZN => n3574);
   U15919 : OAI22_X1 port map( A1 => n18594, A2 => n16669, B1 => n16779, B2 => 
                           n16670, ZN => n3573);
   U15920 : OAI22_X1 port map( A1 => n18595, A2 => n16671, B1 => n16781, B2 => 
                           n16672, ZN => n3572);
   U15921 : OAI22_X1 port map( A1 => n17494, A2 => n16671, B1 => n16782, B2 => 
                           n16672, ZN => n3571);
   U15922 : OAI22_X1 port map( A1 => n17495, A2 => n16669, B1 => n16783, B2 => 
                           n16672, ZN => n3570);
   U15923 : OAI22_X1 port map( A1 => n17496, A2 => n16671, B1 => n16784, B2 => 
                           n16672, ZN => n3569);
   U15924 : OAI22_X1 port map( A1 => n17848, A2 => n16669, B1 => n16785, B2 => 
                           n16672, ZN => n3568);
   U15925 : OAI22_X1 port map( A1 => n17497, A2 => n16671, B1 => n16786, B2 => 
                           n16672, ZN => n3567);
   U15926 : OAI22_X1 port map( A1 => n17498, A2 => n16669, B1 => n16787, B2 => 
                           n16672, ZN => n3566);
   U15927 : OAI22_X1 port map( A1 => n17239, A2 => n16669, B1 => n16788, B2 => 
                           n16672, ZN => n3565);
   U15928 : OAI22_X1 port map( A1 => n17499, A2 => n16669, B1 => n16789, B2 => 
                           n16672, ZN => n3564);
   U15929 : OAI22_X1 port map( A1 => n17500, A2 => n16669, B1 => n16790, B2 => 
                           n16672, ZN => n3563);
   U15930 : OAI22_X1 port map( A1 => n17240, A2 => n16669, B1 => n16791, B2 => 
                           n16672, ZN => n3562);
   U15931 : OAI22_X1 port map( A1 => n17241, A2 => n16669, B1 => n16792, B2 => 
                           n16672, ZN => n3561);
   U15932 : OAI22_X1 port map( A1 => n17849, A2 => n16669, B1 => n16793, B2 => 
                           n16672, ZN => n3560);
   U15933 : OAI22_X1 port map( A1 => n18596, A2 => n16671, B1 => n16794, B2 => 
                           n16672, ZN => n3559);
   U15934 : OAI22_X1 port map( A1 => n18597, A2 => n16671, B1 => n16795, B2 => 
                           n16672, ZN => n3558);
   U15935 : OAI22_X1 port map( A1 => n18196, A2 => n16669, B1 => n16796, B2 => 
                           n16672, ZN => n3557);
   U15936 : OAI22_X1 port map( A1 => n18598, A2 => n16669, B1 => n16797, B2 => 
                           n16672, ZN => n3556);
   U15937 : OAI22_X1 port map( A1 => n18599, A2 => n16671, B1 => n16798, B2 => 
                           n16672, ZN => n3555);
   U15938 : OAI22_X1 port map( A1 => n18600, A2 => n16669, B1 => n16799, B2 => 
                           n16672, ZN => n3554);
   U15939 : OAI22_X1 port map( A1 => n18197, A2 => n16671, B1 => n16800, B2 => 
                           n16672, ZN => n3553);
   U15940 : OAI22_X1 port map( A1 => n18198, A2 => n16669, B1 => n16801, B2 => 
                           n16672, ZN => n3552);
   U15941 : OAI22_X1 port map( A1 => n18199, A2 => n16671, B1 => n16802, B2 => 
                           n16672, ZN => n3551);
   U15942 : OAI22_X1 port map( A1 => n18601, A2 => n16671, B1 => n16803, B2 => 
                           n16672, ZN => n3550);
   U15943 : OAI22_X1 port map( A1 => n18200, A2 => n16669, B1 => n16804, B2 => 
                           n16672, ZN => n3549);
   U15944 : OAI22_X1 port map( A1 => n18602, A2 => n16669, B1 => n16805, B2 => 
                           n16670, ZN => n3548);
   U15945 : OAI22_X1 port map( A1 => n18603, A2 => n16671, B1 => n16806, B2 => 
                           n16672, ZN => n3547);
   U15946 : OAI22_X1 port map( A1 => n18604, A2 => n16669, B1 => n16808, B2 => 
                           n16672, ZN => n3546);
   U15947 : OAI22_X1 port map( A1 => n18201, A2 => n16671, B1 => n16810, B2 => 
                           n16670, ZN => n3545);
   U15948 : OAI22_X1 port map( A1 => n18202, A2 => n16669, B1 => n16812, B2 => 
                           n16672, ZN => n3544);
   U15949 : NAND2_X1 port map( A1 => n16814, A2 => n16673, ZN => n16675);
   U15950 : CLKBUF_X2 port map( A => n16675, Z => n16677);
   U15951 : NAND2_X1 port map( A1 => n13731, A2 => n16677, ZN => n16676);
   U15952 : OAI22_X1 port map( A1 => n17501, A2 => n16676, B1 => n16815, B2 => 
                           n16675, ZN => n3543);
   U15953 : CLKBUF_X2 port map( A => n16676, Z => n16674);
   U15954 : OAI22_X1 port map( A1 => n17850, A2 => n16674, B1 => n16816, B2 => 
                           n16677, ZN => n3542);
   U15955 : OAI22_X1 port map( A1 => n17502, A2 => n16676, B1 => n16817, B2 => 
                           n16675, ZN => n3541);
   U15956 : OAI22_X1 port map( A1 => n17851, A2 => n16674, B1 => n16818, B2 => 
                           n16675, ZN => n3540);
   U15957 : OAI22_X1 port map( A1 => n17503, A2 => n16674, B1 => n16819, B2 => 
                           n16677, ZN => n3539);
   U15958 : OAI22_X1 port map( A1 => n17504, A2 => n16674, B1 => n16820, B2 => 
                           n16675, ZN => n3538);
   U15959 : OAI22_X1 port map( A1 => n17242, A2 => n16674, B1 => n16821, B2 => 
                           n16677, ZN => n3537);
   U15960 : OAI22_X1 port map( A1 => n17243, A2 => n16674, B1 => n16822, B2 => 
                           n16677, ZN => n3536);
   U15961 : OAI22_X1 port map( A1 => n17852, A2 => n16674, B1 => n16823, B2 => 
                           n16677, ZN => n3535);
   U15962 : OAI22_X1 port map( A1 => n17244, A2 => n16674, B1 => n16824, B2 => 
                           n16677, ZN => n3534);
   U15963 : OAI22_X1 port map( A1 => n17505, A2 => n16674, B1 => n16825, B2 => 
                           n16677, ZN => n3533);
   U15964 : OAI22_X1 port map( A1 => n17853, A2 => n16674, B1 => n16826, B2 => 
                           n16675, ZN => n3532);
   U15965 : OAI22_X1 port map( A1 => n18605, A2 => n16676, B1 => n16827, B2 => 
                           n16675, ZN => n3531);
   U15966 : OAI22_X1 port map( A1 => n18203, A2 => n16674, B1 => n16828, B2 => 
                           n16677, ZN => n3530);
   U15967 : OAI22_X1 port map( A1 => n18606, A2 => n16674, B1 => n16829, B2 => 
                           n16675, ZN => n3529);
   U15968 : OAI22_X1 port map( A1 => n18607, A2 => n16676, B1 => n16830, B2 => 
                           n16675, ZN => n3528);
   U15969 : OAI22_X1 port map( A1 => n18608, A2 => n16676, B1 => n16831, B2 => 
                           n16675, ZN => n3527);
   U15970 : OAI22_X1 port map( A1 => n18861, A2 => n16674, B1 => n16832, B2 => 
                           n16677, ZN => n3526);
   U15971 : OAI22_X1 port map( A1 => n18204, A2 => n16674, B1 => n16833, B2 => 
                           n16675, ZN => n3525);
   U15972 : OAI22_X1 port map( A1 => n18205, A2 => n16676, B1 => n16834, B2 => 
                           n16675, ZN => n3524);
   U15973 : OAI22_X1 port map( A1 => n18862, A2 => n16676, B1 => n16835, B2 => 
                           n16677, ZN => n3523);
   U15974 : OAI22_X1 port map( A1 => n18609, A2 => n16674, B1 => n16836, B2 => 
                           n16677, ZN => n3522);
   U15975 : OAI22_X1 port map( A1 => n18610, A2 => n16674, B1 => n16837, B2 => 
                           n16677, ZN => n3521);
   U15976 : OAI22_X1 port map( A1 => n18863, A2 => n16674, B1 => n16838, B2 => 
                           n16675, ZN => n3520);
   U15977 : OAI22_X1 port map( A1 => n18864, A2 => n16674, B1 => n16839, B2 => 
                           n16677, ZN => n3519);
   U15978 : OAI22_X1 port map( A1 => n18206, A2 => n16676, B1 => n16840, B2 => 
                           n16675, ZN => n3518);
   U15979 : OAI22_X1 port map( A1 => n18611, A2 => n16674, B1 => n16841, B2 => 
                           n16675, ZN => n3517);
   U15980 : OAI22_X1 port map( A1 => n18207, A2 => n16676, B1 => n16842, B2 => 
                           n16675, ZN => n3516);
   U15981 : OAI22_X1 port map( A1 => n18208, A2 => n16674, B1 => n16843, B2 => 
                           n16675, ZN => n3515);
   U15982 : OAI22_X1 port map( A1 => n18612, A2 => n16676, B1 => n16844, B2 => 
                           n16675, ZN => n3514);
   U15983 : OAI22_X1 port map( A1 => n18865, A2 => n16674, B1 => n16845, B2 => 
                           n16675, ZN => n3513);
   U15984 : OAI22_X1 port map( A1 => n18866, A2 => n16676, B1 => n16846, B2 => 
                           n16675, ZN => n3512);
   U15985 : OAI22_X1 port map( A1 => n18613, A2 => n16674, B1 => n16847, B2 => 
                           n16675, ZN => n3511);
   U15986 : OAI22_X1 port map( A1 => n18614, A2 => n16676, B1 => n16848, B2 => 
                           n16675, ZN => n3510);
   U15987 : OAI22_X1 port map( A1 => n18615, A2 => n16674, B1 => n16849, B2 => 
                           n16675, ZN => n3509);
   U15988 : OAI22_X1 port map( A1 => n18867, A2 => n16676, B1 => n16850, B2 => 
                           n16677, ZN => n3508);
   U15989 : OAI22_X1 port map( A1 => n17506, A2 => n16676, B1 => n16851, B2 => 
                           n16677, ZN => n3507);
   U15990 : OAI22_X1 port map( A1 => n17507, A2 => n16674, B1 => n16852, B2 => 
                           n16677, ZN => n3506);
   U15991 : OAI22_X1 port map( A1 => n17245, A2 => n16676, B1 => n16853, B2 => 
                           n16677, ZN => n3505);
   U15992 : OAI22_X1 port map( A1 => n17508, A2 => n16674, B1 => n16854, B2 => 
                           n16677, ZN => n3504);
   U15993 : OAI22_X1 port map( A1 => n17509, A2 => n16676, B1 => n16855, B2 => 
                           n16677, ZN => n3503);
   U15994 : OAI22_X1 port map( A1 => n17854, A2 => n16674, B1 => n16856, B2 => 
                           n16677, ZN => n3502);
   U15995 : OAI22_X1 port map( A1 => n17510, A2 => n16674, B1 => n16857, B2 => 
                           n16677, ZN => n3501);
   U15996 : OAI22_X1 port map( A1 => n17246, A2 => n16674, B1 => n16858, B2 => 
                           n16677, ZN => n3500);
   U15997 : OAI22_X1 port map( A1 => n17855, A2 => n16674, B1 => n16859, B2 => 
                           n16677, ZN => n3499);
   U15998 : OAI22_X1 port map( A1 => n17511, A2 => n16674, B1 => n16860, B2 => 
                           n16677, ZN => n3498);
   U15999 : OAI22_X1 port map( A1 => n17512, A2 => n16674, B1 => n16861, B2 => 
                           n16677, ZN => n3497);
   U16000 : OAI22_X1 port map( A1 => n17856, A2 => n16674, B1 => n16862, B2 => 
                           n16677, ZN => n3496);
   U16001 : OAI22_X1 port map( A1 => n18616, A2 => n16676, B1 => n16863, B2 => 
                           n16677, ZN => n3495);
   U16002 : OAI22_X1 port map( A1 => n18209, A2 => n16676, B1 => n16864, B2 => 
                           n16677, ZN => n3494);
   U16003 : OAI22_X1 port map( A1 => n18868, A2 => n16674, B1 => n16865, B2 => 
                           n16677, ZN => n3493);
   U16004 : OAI22_X1 port map( A1 => n18617, A2 => n16674, B1 => n16866, B2 => 
                           n16677, ZN => n3492);
   U16005 : OAI22_X1 port map( A1 => n18210, A2 => n16676, B1 => n16867, B2 => 
                           n16677, ZN => n3491);
   U16006 : OAI22_X1 port map( A1 => n18211, A2 => n16674, B1 => n16868, B2 => 
                           n16677, ZN => n3490);
   U16007 : OAI22_X1 port map( A1 => n18212, A2 => n16676, B1 => n16869, B2 => 
                           n16677, ZN => n3489);
   U16008 : OAI22_X1 port map( A1 => n18618, A2 => n16674, B1 => n16870, B2 => 
                           n16677, ZN => n3488);
   U16009 : OAI22_X1 port map( A1 => n18213, A2 => n16676, B1 => n16871, B2 => 
                           n16677, ZN => n3487);
   U16010 : OAI22_X1 port map( A1 => n18869, A2 => n16676, B1 => n16872, B2 => 
                           n16677, ZN => n3486);
   U16011 : OAI22_X1 port map( A1 => n18619, A2 => n16674, B1 => n16873, B2 => 
                           n16677, ZN => n3485);
   U16012 : OAI22_X1 port map( A1 => n18870, A2 => n16674, B1 => n16874, B2 => 
                           n16675, ZN => n3484);
   U16013 : OAI22_X1 port map( A1 => n18620, A2 => n16676, B1 => n16875, B2 => 
                           n16677, ZN => n3483);
   U16014 : OAI22_X1 port map( A1 => n18871, A2 => n16674, B1 => n16876, B2 => 
                           n16677, ZN => n3482);
   U16015 : OAI22_X1 port map( A1 => n18621, A2 => n16676, B1 => n16878, B2 => 
                           n16675, ZN => n3481);
   U16016 : OAI22_X1 port map( A1 => n18622, A2 => n16674, B1 => n16881, B2 => 
                           n16677, ZN => n3480);
   U16017 : NAND2_X1 port map( A1 => WR, A2 => ADD_WR(4), ZN => n16712);
   U16018 : NAND2_X1 port map( A1 => n16714, A2 => n16707, ZN => n16680);
   U16019 : CLKBUF_X2 port map( A => n16680, Z => n16682);
   U16020 : NAND2_X1 port map( A1 => n13731, A2 => n16682, ZN => n16681);
   U16021 : OAI22_X1 port map( A1 => n17513, A2 => n16681, B1 => n16815, B2 => 
                           n16680, ZN => n3479);
   U16022 : CLKBUF_X2 port map( A => n16681, Z => n16679);
   U16023 : OAI22_X1 port map( A1 => n17514, A2 => n16679, B1 => n16816, B2 => 
                           n16682, ZN => n3478);
   U16024 : OAI22_X1 port map( A1 => n17515, A2 => n16681, B1 => n16817, B2 => 
                           n16680, ZN => n3477);
   U16025 : OAI22_X1 port map( A1 => n17247, A2 => n16679, B1 => n16818, B2 => 
                           n16680, ZN => n3476);
   U16026 : OAI22_X1 port map( A1 => n17248, A2 => n16679, B1 => n16819, B2 => 
                           n16682, ZN => n3475);
   U16027 : OAI22_X1 port map( A1 => n17516, A2 => n16679, B1 => n16820, B2 => 
                           n16680, ZN => n3474);
   U16028 : OAI22_X1 port map( A1 => n17517, A2 => n16679, B1 => n16821, B2 => 
                           n16682, ZN => n3473);
   U16029 : OAI22_X1 port map( A1 => n17857, A2 => n16679, B1 => n16822, B2 => 
                           n16682, ZN => n3472);
   U16030 : OAI22_X1 port map( A1 => n17518, A2 => n16679, B1 => n16823, B2 => 
                           n16682, ZN => n3471);
   U16031 : OAI22_X1 port map( A1 => n17858, A2 => n16679, B1 => n16824, B2 => 
                           n16682, ZN => n3470);
   U16032 : OAI22_X1 port map( A1 => n17519, A2 => n16679, B1 => n16825, B2 => 
                           n16682, ZN => n3469);
   U16033 : OAI22_X1 port map( A1 => n17520, A2 => n16679, B1 => n16826, B2 => 
                           n16680, ZN => n3468);
   U16034 : OAI22_X1 port map( A1 => n18214, A2 => n16681, B1 => n16827, B2 => 
                           n16680, ZN => n3467);
   U16035 : OAI22_X1 port map( A1 => n18215, A2 => n16679, B1 => n16828, B2 => 
                           n16682, ZN => n3466);
   U16036 : OAI22_X1 port map( A1 => n18623, A2 => n16679, B1 => n16829, B2 => 
                           n16680, ZN => n3465);
   U16037 : OAI22_X1 port map( A1 => n18216, A2 => n16681, B1 => n16830, B2 => 
                           n16680, ZN => n3464);
   U16038 : OAI22_X1 port map( A1 => n18624, A2 => n16681, B1 => n16831, B2 => 
                           n16680, ZN => n3463);
   U16039 : OAI22_X1 port map( A1 => n18625, A2 => n16679, B1 => n16832, B2 => 
                           n16682, ZN => n3462);
   U16040 : OAI22_X1 port map( A1 => n18872, A2 => n16679, B1 => n16833, B2 => 
                           n16680, ZN => n3461);
   U16041 : OAI22_X1 port map( A1 => n18217, A2 => n16681, B1 => n16834, B2 => 
                           n16680, ZN => n3460);
   U16042 : OAI22_X1 port map( A1 => n18626, A2 => n16681, B1 => n16835, B2 => 
                           n16682, ZN => n3459);
   U16043 : OAI22_X1 port map( A1 => n18627, A2 => n16679, B1 => n16836, B2 => 
                           n16682, ZN => n3458);
   U16044 : OAI22_X1 port map( A1 => n18628, A2 => n16679, B1 => n16837, B2 => 
                           n16682, ZN => n3457);
   U16045 : OAI22_X1 port map( A1 => n18218, A2 => n16679, B1 => n16838, B2 => 
                           n16680, ZN => n3456);
   U16046 : OAI22_X1 port map( A1 => n18219, A2 => n16679, B1 => n16839, B2 => 
                           n16682, ZN => n3455);
   U16047 : OAI22_X1 port map( A1 => n18629, A2 => n16681, B1 => n16840, B2 => 
                           n16680, ZN => n3454);
   U16048 : OAI22_X1 port map( A1 => n18873, A2 => n16679, B1 => n16841, B2 => 
                           n16680, ZN => n3453);
   U16049 : OAI22_X1 port map( A1 => n18630, A2 => n16681, B1 => n16842, B2 => 
                           n16680, ZN => n3452);
   U16050 : OAI22_X1 port map( A1 => n18220, A2 => n16679, B1 => n16843, B2 => 
                           n16680, ZN => n3451);
   U16051 : OAI22_X1 port map( A1 => n18221, A2 => n16681, B1 => n16844, B2 => 
                           n16680, ZN => n3450);
   U16052 : OAI22_X1 port map( A1 => n18631, A2 => n16679, B1 => n16845, B2 => 
                           n16680, ZN => n3449);
   U16053 : OAI22_X1 port map( A1 => n18632, A2 => n16681, B1 => n16846, B2 => 
                           n16680, ZN => n3448);
   U16054 : OAI22_X1 port map( A1 => n18874, A2 => n16679, B1 => n16847, B2 => 
                           n16680, ZN => n3447);
   U16055 : OAI22_X1 port map( A1 => n18633, A2 => n16681, B1 => n16848, B2 => 
                           n16680, ZN => n3446);
   U16056 : OAI22_X1 port map( A1 => n18222, A2 => n16679, B1 => n16849, B2 => 
                           n16680, ZN => n3445);
   U16057 : OAI22_X1 port map( A1 => n18634, A2 => n16681, B1 => n16850, B2 => 
                           n16682, ZN => n3444);
   U16058 : OAI22_X1 port map( A1 => n17249, A2 => n16681, B1 => n16851, B2 => 
                           n16682, ZN => n3443);
   U16059 : OAI22_X1 port map( A1 => n17859, A2 => n16679, B1 => n16852, B2 => 
                           n16682, ZN => n3442);
   U16060 : OAI22_X1 port map( A1 => n17521, A2 => n16681, B1 => n16853, B2 => 
                           n16682, ZN => n3441);
   U16061 : OAI22_X1 port map( A1 => n17522, A2 => n16679, B1 => n16854, B2 => 
                           n16682, ZN => n3440);
   U16062 : OAI22_X1 port map( A1 => n17860, A2 => n16681, B1 => n16855, B2 => 
                           n16682, ZN => n3439);
   U16063 : OAI22_X1 port map( A1 => n17861, A2 => n16679, B1 => n16856, B2 => 
                           n16682, ZN => n3438);
   U16064 : OAI22_X1 port map( A1 => n17523, A2 => n16679, B1 => n16857, B2 => 
                           n16682, ZN => n3437);
   U16065 : OAI22_X1 port map( A1 => n17524, A2 => n16679, B1 => n16858, B2 => 
                           n16682, ZN => n3436);
   U16066 : OAI22_X1 port map( A1 => n17525, A2 => n16679, B1 => n16859, B2 => 
                           n16682, ZN => n3435);
   U16067 : OAI22_X1 port map( A1 => n17526, A2 => n16679, B1 => n16860, B2 => 
                           n16682, ZN => n3434);
   U16068 : OAI22_X1 port map( A1 => n17527, A2 => n16679, B1 => n16861, B2 => 
                           n16682, ZN => n3433);
   U16069 : OAI22_X1 port map( A1 => n17250, A2 => n16679, B1 => n16862, B2 => 
                           n16682, ZN => n3432);
   U16070 : OAI22_X1 port map( A1 => n18223, A2 => n16681, B1 => n16863, B2 => 
                           n16682, ZN => n3431);
   U16071 : OAI22_X1 port map( A1 => n18635, A2 => n16681, B1 => n16864, B2 => 
                           n16682, ZN => n3430);
   U16072 : OAI22_X1 port map( A1 => n18224, A2 => n16679, B1 => n16865, B2 => 
                           n16682, ZN => n3429);
   U16073 : OAI22_X1 port map( A1 => n18225, A2 => n16679, B1 => n16866, B2 => 
                           n16682, ZN => n3428);
   U16074 : OAI22_X1 port map( A1 => n18636, A2 => n16681, B1 => n16867, B2 => 
                           n16682, ZN => n3427);
   U16075 : OAI22_X1 port map( A1 => n18637, A2 => n16679, B1 => n16868, B2 => 
                           n16682, ZN => n3426);
   U16076 : OAI22_X1 port map( A1 => n18875, A2 => n16681, B1 => n16869, B2 => 
                           n16682, ZN => n3425);
   U16077 : OAI22_X1 port map( A1 => n18876, A2 => n16679, B1 => n16870, B2 => 
                           n16682, ZN => n3424);
   U16078 : OAI22_X1 port map( A1 => n18226, A2 => n16681, B1 => n16871, B2 => 
                           n16682, ZN => n3423);
   U16079 : OAI22_X1 port map( A1 => n18227, A2 => n16681, B1 => n16872, B2 => 
                           n16682, ZN => n3422);
   U16080 : OAI22_X1 port map( A1 => n18228, A2 => n16679, B1 => n16873, B2 => 
                           n16682, ZN => n3421);
   U16081 : OAI22_X1 port map( A1 => n18638, A2 => n16679, B1 => n16874, B2 => 
                           n16680, ZN => n3420);
   U16082 : OAI22_X1 port map( A1 => n18639, A2 => n16681, B1 => n16875, B2 => 
                           n16682, ZN => n3419);
   U16083 : OAI22_X1 port map( A1 => n18640, A2 => n16679, B1 => n16876, B2 => 
                           n16682, ZN => n3418);
   U16084 : OAI22_X1 port map( A1 => n18641, A2 => n16681, B1 => n16878, B2 => 
                           n16680, ZN => n3417);
   U16085 : OAI22_X1 port map( A1 => n18229, A2 => n16679, B1 => n16881, B2 => 
                           n16682, ZN => n3416);
   U16086 : NAND2_X1 port map( A1 => n16719, A2 => n16707, ZN => n16684);
   U16087 : CLKBUF_X2 port map( A => n16684, Z => n16686);
   U16088 : NAND2_X1 port map( A1 => n13731, A2 => n16686, ZN => n16685);
   U16089 : OAI22_X1 port map( A1 => n17251, A2 => n16685, B1 => n16745, B2 => 
                           n16684, ZN => n3415);
   U16090 : CLKBUF_X2 port map( A => n16685, Z => n16683);
   U16091 : OAI22_X1 port map( A1 => n17862, A2 => n16683, B1 => n16746, B2 => 
                           n16686, ZN => n3414);
   U16092 : OAI22_X1 port map( A1 => n17528, A2 => n16685, B1 => n16747, B2 => 
                           n16684, ZN => n3413);
   U16093 : OAI22_X1 port map( A1 => n17529, A2 => n16683, B1 => n16748, B2 => 
                           n16684, ZN => n3412);
   U16094 : OAI22_X1 port map( A1 => n17530, A2 => n16683, B1 => n16749, B2 => 
                           n16686, ZN => n3411);
   U16095 : OAI22_X1 port map( A1 => n17531, A2 => n16683, B1 => n16750, B2 => 
                           n16684, ZN => n3410);
   U16096 : OAI22_X1 port map( A1 => n17863, A2 => n16683, B1 => n16751, B2 => 
                           n16686, ZN => n3409);
   U16097 : OAI22_X1 port map( A1 => n17864, A2 => n16683, B1 => n16752, B2 => 
                           n16686, ZN => n3408);
   U16098 : OAI22_X1 port map( A1 => n17532, A2 => n16683, B1 => n16753, B2 => 
                           n16686, ZN => n3407);
   U16099 : OAI22_X1 port map( A1 => n17865, A2 => n16683, B1 => n16754, B2 => 
                           n16686, ZN => n3406);
   U16100 : OAI22_X1 port map( A1 => n17533, A2 => n16683, B1 => n16755, B2 => 
                           n16686, ZN => n3405);
   U16101 : OAI22_X1 port map( A1 => n17866, A2 => n16683, B1 => n16756, B2 => 
                           n16684, ZN => n3404);
   U16102 : OAI22_X1 port map( A1 => n18877, A2 => n16685, B1 => n16757, B2 => 
                           n16684, ZN => n3403);
   U16103 : OAI22_X1 port map( A1 => n18878, A2 => n16683, B1 => n16758, B2 => 
                           n16686, ZN => n3402);
   U16104 : OAI22_X1 port map( A1 => n18879, A2 => n16683, B1 => n16759, B2 => 
                           n16684, ZN => n3401);
   U16105 : OAI22_X1 port map( A1 => n18880, A2 => n16685, B1 => n16760, B2 => 
                           n16684, ZN => n3400);
   U16106 : OAI22_X1 port map( A1 => n18881, A2 => n16685, B1 => n16761, B2 => 
                           n16684, ZN => n3399);
   U16107 : OAI22_X1 port map( A1 => n18882, A2 => n16683, B1 => n16762, B2 => 
                           n16686, ZN => n3398);
   U16108 : OAI22_X1 port map( A1 => n18883, A2 => n16683, B1 => n16763, B2 => 
                           n16684, ZN => n3397);
   U16109 : OAI22_X1 port map( A1 => n18884, A2 => n16685, B1 => n16764, B2 => 
                           n16684, ZN => n3396);
   U16110 : OAI22_X1 port map( A1 => n18885, A2 => n16685, B1 => n16765, B2 => 
                           n16686, ZN => n3395);
   U16111 : OAI22_X1 port map( A1 => n18642, A2 => n16683, B1 => n16766, B2 => 
                           n16686, ZN => n3394);
   U16112 : OAI22_X1 port map( A1 => n18643, A2 => n16683, B1 => n16767, B2 => 
                           n16686, ZN => n3393);
   U16113 : OAI22_X1 port map( A1 => n18644, A2 => n16683, B1 => n16768, B2 => 
                           n16684, ZN => n3392);
   U16114 : OAI22_X1 port map( A1 => n18645, A2 => n16683, B1 => n16769, B2 => 
                           n16686, ZN => n3391);
   U16115 : OAI22_X1 port map( A1 => n18646, A2 => n16685, B1 => n16770, B2 => 
                           n16684, ZN => n3390);
   U16116 : OAI22_X1 port map( A1 => n18886, A2 => n16683, B1 => n16771, B2 => 
                           n16684, ZN => n3389);
   U16117 : OAI22_X1 port map( A1 => n18647, A2 => n16685, B1 => n16772, B2 => 
                           n16684, ZN => n3388);
   U16118 : OAI22_X1 port map( A1 => n18648, A2 => n16683, B1 => n16773, B2 => 
                           n16684, ZN => n3387);
   U16119 : OAI22_X1 port map( A1 => n18649, A2 => n16685, B1 => n16774, B2 => 
                           n16684, ZN => n3386);
   U16120 : OAI22_X1 port map( A1 => n18650, A2 => n16683, B1 => n16775, B2 => 
                           n16684, ZN => n3385);
   U16121 : OAI22_X1 port map( A1 => n18887, A2 => n16685, B1 => n16776, B2 => 
                           n16684, ZN => n3384);
   U16122 : OAI22_X1 port map( A1 => n18651, A2 => n16683, B1 => n16777, B2 => 
                           n16684, ZN => n3383);
   U16123 : OAI22_X1 port map( A1 => n18888, A2 => n16685, B1 => n16778, B2 => 
                           n16684, ZN => n3382);
   U16124 : OAI22_X1 port map( A1 => n18889, A2 => n16683, B1 => n16779, B2 => 
                           n16684, ZN => n3381);
   U16125 : OAI22_X1 port map( A1 => n18890, A2 => n16685, B1 => n16781, B2 => 
                           n16686, ZN => n3380);
   U16126 : OAI22_X1 port map( A1 => n17534, A2 => n16685, B1 => n16782, B2 => 
                           n16686, ZN => n3379);
   U16127 : OAI22_X1 port map( A1 => n17252, A2 => n16683, B1 => n16783, B2 => 
                           n16686, ZN => n3378);
   U16128 : OAI22_X1 port map( A1 => n17535, A2 => n16685, B1 => n16784, B2 => 
                           n16686, ZN => n3377);
   U16129 : OAI22_X1 port map( A1 => n17253, A2 => n16683, B1 => n16785, B2 => 
                           n16686, ZN => n3376);
   U16130 : OAI22_X1 port map( A1 => n17867, A2 => n16685, B1 => n16786, B2 => 
                           n16686, ZN => n3375);
   U16131 : OAI22_X1 port map( A1 => n17536, A2 => n16683, B1 => n16787, B2 => 
                           n16686, ZN => n3374);
   U16132 : OAI22_X1 port map( A1 => n17537, A2 => n16683, B1 => n16788, B2 => 
                           n16686, ZN => n3373);
   U16133 : OAI22_X1 port map( A1 => n17538, A2 => n16683, B1 => n16789, B2 => 
                           n16686, ZN => n3372);
   U16134 : OAI22_X1 port map( A1 => n17868, A2 => n16683, B1 => n16790, B2 => 
                           n16686, ZN => n3371);
   U16135 : OAI22_X1 port map( A1 => n17539, A2 => n16683, B1 => n16791, B2 => 
                           n16686, ZN => n3370);
   U16136 : OAI22_X1 port map( A1 => n17869, A2 => n16683, B1 => n16792, B2 => 
                           n16686, ZN => n3369);
   U16137 : OAI22_X1 port map( A1 => n17540, A2 => n16683, B1 => n16793, B2 => 
                           n16686, ZN => n3368);
   U16138 : OAI22_X1 port map( A1 => n18652, A2 => n16685, B1 => n16794, B2 => 
                           n16686, ZN => n3367);
   U16139 : OAI22_X1 port map( A1 => n18653, A2 => n16685, B1 => n16795, B2 => 
                           n16686, ZN => n3366);
   U16140 : OAI22_X1 port map( A1 => n18891, A2 => n16683, B1 => n16796, B2 => 
                           n16686, ZN => n3365);
   U16141 : OAI22_X1 port map( A1 => n18654, A2 => n16683, B1 => n16797, B2 => 
                           n16686, ZN => n3364);
   U16142 : OAI22_X1 port map( A1 => n18892, A2 => n16685, B1 => n16798, B2 => 
                           n16686, ZN => n3363);
   U16143 : OAI22_X1 port map( A1 => n18893, A2 => n16683, B1 => n16799, B2 => 
                           n16686, ZN => n3362);
   U16144 : OAI22_X1 port map( A1 => n18655, A2 => n16685, B1 => n16800, B2 => 
                           n16686, ZN => n3361);
   U16145 : OAI22_X1 port map( A1 => n18656, A2 => n16683, B1 => n16801, B2 => 
                           n16686, ZN => n3360);
   U16146 : OAI22_X1 port map( A1 => n18894, A2 => n16685, B1 => n16802, B2 => 
                           n16686, ZN => n3359);
   U16147 : OAI22_X1 port map( A1 => n18895, A2 => n16685, B1 => n16803, B2 => 
                           n16686, ZN => n3358);
   U16148 : OAI22_X1 port map( A1 => n18230, A2 => n16683, B1 => n16804, B2 => 
                           n16686, ZN => n3357);
   U16149 : OAI22_X1 port map( A1 => n18896, A2 => n16683, B1 => n16805, B2 => 
                           n16684, ZN => n3356);
   U16150 : OAI22_X1 port map( A1 => n18657, A2 => n16685, B1 => n16806, B2 => 
                           n16686, ZN => n3355);
   U16151 : OAI22_X1 port map( A1 => n18658, A2 => n16683, B1 => n16808, B2 => 
                           n16686, ZN => n3354);
   U16152 : OAI22_X1 port map( A1 => n18659, A2 => n16685, B1 => n16810, B2 => 
                           n16684, ZN => n3353);
   U16153 : OAI22_X1 port map( A1 => n18897, A2 => n16683, B1 => n16812, B2 => 
                           n16686, ZN => n3352);
   U16154 : NAND2_X1 port map( A1 => n16724, A2 => n16707, ZN => n16688);
   U16155 : CLKBUF_X2 port map( A => n16688, Z => n16690);
   U16156 : NAND2_X1 port map( A1 => n13731, A2 => n16690, ZN => n16689);
   U16157 : OAI22_X1 port map( A1 => n17541, A2 => n16689, B1 => n16745, B2 => 
                           n16688, ZN => n3351);
   U16158 : CLKBUF_X2 port map( A => n16689, Z => n16687);
   U16159 : OAI22_X1 port map( A1 => n17870, A2 => n16687, B1 => n16746, B2 => 
                           n16690, ZN => n3350);
   U16160 : OAI22_X1 port map( A1 => n17542, A2 => n16689, B1 => n16747, B2 => 
                           n16688, ZN => n3349);
   U16161 : OAI22_X1 port map( A1 => n17543, A2 => n16687, B1 => n16748, B2 => 
                           n16688, ZN => n3348);
   U16162 : OAI22_X1 port map( A1 => n17254, A2 => n16687, B1 => n16749, B2 => 
                           n16690, ZN => n3347);
   U16163 : OAI22_X1 port map( A1 => n17544, A2 => n16687, B1 => n16750, B2 => 
                           n16688, ZN => n3346);
   U16164 : OAI22_X1 port map( A1 => n17871, A2 => n16687, B1 => n16751, B2 => 
                           n16690, ZN => n3345);
   U16165 : OAI22_X1 port map( A1 => n17255, A2 => n16687, B1 => n16752, B2 => 
                           n16690, ZN => n3344);
   U16166 : OAI22_X1 port map( A1 => n17545, A2 => n16687, B1 => n16753, B2 => 
                           n16690, ZN => n3343);
   U16167 : OAI22_X1 port map( A1 => n17872, A2 => n16687, B1 => n16754, B2 => 
                           n16690, ZN => n3342);
   U16168 : OAI22_X1 port map( A1 => n17546, A2 => n16687, B1 => n16755, B2 => 
                           n16690, ZN => n3341);
   U16169 : OAI22_X1 port map( A1 => n17873, A2 => n16687, B1 => n16756, B2 => 
                           n16688, ZN => n3340);
   U16170 : OAI22_X1 port map( A1 => n18898, A2 => n16689, B1 => n16757, B2 => 
                           n16688, ZN => n3339);
   U16171 : OAI22_X1 port map( A1 => n18660, A2 => n16687, B1 => n16758, B2 => 
                           n16690, ZN => n3338);
   U16172 : OAI22_X1 port map( A1 => n18661, A2 => n16687, B1 => n16759, B2 => 
                           n16688, ZN => n3337);
   U16173 : OAI22_X1 port map( A1 => n18231, A2 => n16689, B1 => n16760, B2 => 
                           n16688, ZN => n3336);
   U16174 : OAI22_X1 port map( A1 => n18662, A2 => n16689, B1 => n16761, B2 => 
                           n16688, ZN => n3335);
   U16175 : OAI22_X1 port map( A1 => n18899, A2 => n16687, B1 => n16762, B2 => 
                           n16690, ZN => n3334);
   U16176 : OAI22_X1 port map( A1 => n18900, A2 => n16687, B1 => n16763, B2 => 
                           n16688, ZN => n3333);
   U16177 : OAI22_X1 port map( A1 => n18901, A2 => n16689, B1 => n16764, B2 => 
                           n16688, ZN => n3332);
   U16178 : OAI22_X1 port map( A1 => n18902, A2 => n16689, B1 => n16765, B2 => 
                           n16690, ZN => n3331);
   U16179 : OAI22_X1 port map( A1 => n18663, A2 => n16687, B1 => n16766, B2 => 
                           n16690, ZN => n3330);
   U16180 : OAI22_X1 port map( A1 => n18903, A2 => n16687, B1 => n16767, B2 => 
                           n16690, ZN => n3329);
   U16181 : OAI22_X1 port map( A1 => n18664, A2 => n16687, B1 => n16768, B2 => 
                           n16688, ZN => n3328);
   U16182 : OAI22_X1 port map( A1 => n18904, A2 => n16687, B1 => n16769, B2 => 
                           n16690, ZN => n3327);
   U16183 : OAI22_X1 port map( A1 => n18905, A2 => n16689, B1 => n16770, B2 => 
                           n16688, ZN => n3326);
   U16184 : OAI22_X1 port map( A1 => n18665, A2 => n16687, B1 => n16771, B2 => 
                           n16688, ZN => n3325);
   U16185 : OAI22_X1 port map( A1 => n18906, A2 => n16689, B1 => n16772, B2 => 
                           n16688, ZN => n3324);
   U16186 : OAI22_X1 port map( A1 => n18666, A2 => n16687, B1 => n16773, B2 => 
                           n16688, ZN => n3323);
   U16187 : OAI22_X1 port map( A1 => n18667, A2 => n16689, B1 => n16774, B2 => 
                           n16688, ZN => n3322);
   U16188 : OAI22_X1 port map( A1 => n18232, A2 => n16687, B1 => n16775, B2 => 
                           n16688, ZN => n3321);
   U16189 : OAI22_X1 port map( A1 => n18907, A2 => n16689, B1 => n16776, B2 => 
                           n16688, ZN => n3320);
   U16190 : OAI22_X1 port map( A1 => n18668, A2 => n16687, B1 => n16777, B2 => 
                           n16688, ZN => n3319);
   U16191 : OAI22_X1 port map( A1 => n18908, A2 => n16689, B1 => n16778, B2 => 
                           n16688, ZN => n3318);
   U16192 : OAI22_X1 port map( A1 => n18909, A2 => n16687, B1 => n16779, B2 => 
                           n16688, ZN => n3317);
   U16193 : OAI22_X1 port map( A1 => n18910, A2 => n16689, B1 => n16781, B2 => 
                           n16690, ZN => n3316);
   U16194 : OAI22_X1 port map( A1 => n17547, A2 => n16689, B1 => n16782, B2 => 
                           n16690, ZN => n3315);
   U16195 : OAI22_X1 port map( A1 => n17548, A2 => n16687, B1 => n16783, B2 => 
                           n16690, ZN => n3314);
   U16196 : OAI22_X1 port map( A1 => n17874, A2 => n16689, B1 => n16784, B2 => 
                           n16690, ZN => n3313);
   U16197 : OAI22_X1 port map( A1 => n17875, A2 => n16687, B1 => n16785, B2 => 
                           n16690, ZN => n3312);
   U16198 : OAI22_X1 port map( A1 => n17549, A2 => n16689, B1 => n16786, B2 => 
                           n16690, ZN => n3311);
   U16199 : OAI22_X1 port map( A1 => n17550, A2 => n16687, B1 => n16787, B2 => 
                           n16690, ZN => n3310);
   U16200 : OAI22_X1 port map( A1 => n17551, A2 => n16687, B1 => n16788, B2 => 
                           n16690, ZN => n3309);
   U16201 : OAI22_X1 port map( A1 => n17876, A2 => n16687, B1 => n16789, B2 => 
                           n16690, ZN => n3308);
   U16202 : OAI22_X1 port map( A1 => n17552, A2 => n16687, B1 => n16790, B2 => 
                           n16690, ZN => n3307);
   U16203 : OAI22_X1 port map( A1 => n17553, A2 => n16687, B1 => n16791, B2 => 
                           n16690, ZN => n3306);
   U16204 : OAI22_X1 port map( A1 => n17554, A2 => n16687, B1 => n16792, B2 => 
                           n16690, ZN => n3305);
   U16205 : OAI22_X1 port map( A1 => n17877, A2 => n16687, B1 => n16793, B2 => 
                           n16690, ZN => n3304);
   U16206 : OAI22_X1 port map( A1 => n18669, A2 => n16689, B1 => n16794, B2 => 
                           n16690, ZN => n3303);
   U16207 : OAI22_X1 port map( A1 => n18670, A2 => n16689, B1 => n16795, B2 => 
                           n16690, ZN => n3302);
   U16208 : OAI22_X1 port map( A1 => n18911, A2 => n16687, B1 => n16796, B2 => 
                           n16690, ZN => n3301);
   U16209 : OAI22_X1 port map( A1 => n18671, A2 => n16687, B1 => n16797, B2 => 
                           n16690, ZN => n3300);
   U16210 : OAI22_X1 port map( A1 => n18912, A2 => n16689, B1 => n16798, B2 => 
                           n16690, ZN => n3299);
   U16211 : OAI22_X1 port map( A1 => n18672, A2 => n16687, B1 => n16799, B2 => 
                           n16690, ZN => n3298);
   U16212 : OAI22_X1 port map( A1 => n18913, A2 => n16689, B1 => n16800, B2 => 
                           n16690, ZN => n3297);
   U16213 : OAI22_X1 port map( A1 => n18673, A2 => n16687, B1 => n16801, B2 => 
                           n16690, ZN => n3296);
   U16214 : OAI22_X1 port map( A1 => n18674, A2 => n16689, B1 => n16802, B2 => 
                           n16690, ZN => n3295);
   U16215 : OAI22_X1 port map( A1 => n18675, A2 => n16689, B1 => n16803, B2 => 
                           n16690, ZN => n3294);
   U16216 : OAI22_X1 port map( A1 => n18676, A2 => n16687, B1 => n16804, B2 => 
                           n16690, ZN => n3293);
   U16217 : OAI22_X1 port map( A1 => n18677, A2 => n16687, B1 => n16805, B2 => 
                           n16688, ZN => n3292);
   U16218 : OAI22_X1 port map( A1 => n18914, A2 => n16689, B1 => n16806, B2 => 
                           n16690, ZN => n3291);
   U16219 : OAI22_X1 port map( A1 => n18915, A2 => n16687, B1 => n16808, B2 => 
                           n16690, ZN => n3290);
   U16220 : OAI22_X1 port map( A1 => n18678, A2 => n16689, B1 => n16810, B2 => 
                           n16688, ZN => n3289);
   U16221 : OAI22_X1 port map( A1 => n18916, A2 => n16687, B1 => n16812, B2 => 
                           n16690, ZN => n3288);
   U16222 : NAND2_X1 port map( A1 => n16729, A2 => n16707, ZN => n16692);
   U16223 : CLKBUF_X2 port map( A => n16692, Z => n16694);
   U16224 : NAND2_X1 port map( A1 => n13731, A2 => n16694, ZN => n16693);
   U16225 : OAI22_X1 port map( A1 => n17555, A2 => n16693, B1 => n16745, B2 => 
                           n16692, ZN => n3287);
   U16226 : CLKBUF_X2 port map( A => n16693, Z => n16691);
   U16227 : OAI22_X1 port map( A1 => n17556, A2 => n16691, B1 => n16746, B2 => 
                           n16694, ZN => n3286);
   U16228 : OAI22_X1 port map( A1 => n17878, A2 => n16693, B1 => n16747, B2 => 
                           n16692, ZN => n3285);
   U16229 : OAI22_X1 port map( A1 => n17557, A2 => n16691, B1 => n16748, B2 => 
                           n16692, ZN => n3284);
   U16230 : OAI22_X1 port map( A1 => n17558, A2 => n16691, B1 => n16749, B2 => 
                           n16694, ZN => n3283);
   U16231 : OAI22_X1 port map( A1 => n17879, A2 => n16691, B1 => n16750, B2 => 
                           n16692, ZN => n3282);
   U16232 : OAI22_X1 port map( A1 => n17880, A2 => n16691, B1 => n16751, B2 => 
                           n16694, ZN => n3281);
   U16233 : OAI22_X1 port map( A1 => n17881, A2 => n16691, B1 => n16752, B2 => 
                           n16694, ZN => n3280);
   U16234 : OAI22_X1 port map( A1 => n17559, A2 => n16691, B1 => n16753, B2 => 
                           n16694, ZN => n3279);
   U16235 : OAI22_X1 port map( A1 => n17882, A2 => n16691, B1 => n16754, B2 => 
                           n16694, ZN => n3278);
   U16236 : OAI22_X1 port map( A1 => n17560, A2 => n16691, B1 => n16755, B2 => 
                           n16694, ZN => n3277);
   U16237 : OAI22_X1 port map( A1 => n17561, A2 => n16691, B1 => n16756, B2 => 
                           n16692, ZN => n3276);
   U16238 : OAI22_X1 port map( A1 => n18917, A2 => n16693, B1 => n16757, B2 => 
                           n16692, ZN => n3275);
   U16239 : OAI22_X1 port map( A1 => n18679, A2 => n16691, B1 => n16758, B2 => 
                           n16694, ZN => n3274);
   U16240 : OAI22_X1 port map( A1 => n18233, A2 => n16691, B1 => n16759, B2 => 
                           n16692, ZN => n3273);
   U16241 : OAI22_X1 port map( A1 => n18680, A2 => n16693, B1 => n16760, B2 => 
                           n16692, ZN => n3272);
   U16242 : OAI22_X1 port map( A1 => n18918, A2 => n16693, B1 => n16761, B2 => 
                           n16692, ZN => n3271);
   U16243 : OAI22_X1 port map( A1 => n18681, A2 => n16691, B1 => n16762, B2 => 
                           n16694, ZN => n3270);
   U16244 : OAI22_X1 port map( A1 => n18682, A2 => n16691, B1 => n16763, B2 => 
                           n16692, ZN => n3269);
   U16245 : OAI22_X1 port map( A1 => n18683, A2 => n16693, B1 => n16764, B2 => 
                           n16692, ZN => n3268);
   U16246 : OAI22_X1 port map( A1 => n18919, A2 => n16693, B1 => n16765, B2 => 
                           n16694, ZN => n3267);
   U16247 : OAI22_X1 port map( A1 => n18920, A2 => n16691, B1 => n16766, B2 => 
                           n16694, ZN => n3266);
   U16248 : OAI22_X1 port map( A1 => n18234, A2 => n16691, B1 => n16767, B2 => 
                           n16694, ZN => n3265);
   U16249 : OAI22_X1 port map( A1 => n18235, A2 => n16691, B1 => n16768, B2 => 
                           n16692, ZN => n3264);
   U16250 : OAI22_X1 port map( A1 => n18921, A2 => n16691, B1 => n16769, B2 => 
                           n16694, ZN => n3263);
   U16251 : OAI22_X1 port map( A1 => n18684, A2 => n16693, B1 => n16770, B2 => 
                           n16692, ZN => n3262);
   U16252 : OAI22_X1 port map( A1 => n18922, A2 => n16691, B1 => n16771, B2 => 
                           n16692, ZN => n3261);
   U16253 : OAI22_X1 port map( A1 => n18923, A2 => n16693, B1 => n16772, B2 => 
                           n16692, ZN => n3260);
   U16254 : OAI22_X1 port map( A1 => n18236, A2 => n16691, B1 => n16773, B2 => 
                           n16692, ZN => n3259);
   U16255 : OAI22_X1 port map( A1 => n18685, A2 => n16693, B1 => n16774, B2 => 
                           n16692, ZN => n3258);
   U16256 : OAI22_X1 port map( A1 => n18686, A2 => n16691, B1 => n16775, B2 => 
                           n16692, ZN => n3257);
   U16257 : OAI22_X1 port map( A1 => n18687, A2 => n16693, B1 => n16776, B2 => 
                           n16692, ZN => n3256);
   U16258 : OAI22_X1 port map( A1 => n18924, A2 => n16691, B1 => n16777, B2 => 
                           n16692, ZN => n3255);
   U16259 : OAI22_X1 port map( A1 => n18237, A2 => n16693, B1 => n16778, B2 => 
                           n16692, ZN => n3254);
   U16260 : OAI22_X1 port map( A1 => n18688, A2 => n16691, B1 => n16779, B2 => 
                           n16692, ZN => n3253);
   U16261 : OAI22_X1 port map( A1 => n18689, A2 => n16693, B1 => n16781, B2 => 
                           n16694, ZN => n3252);
   U16262 : OAI22_X1 port map( A1 => n17883, A2 => n16693, B1 => n16782, B2 => 
                           n16694, ZN => n3251);
   U16263 : OAI22_X1 port map( A1 => n17562, A2 => n16691, B1 => n16783, B2 => 
                           n16694, ZN => n3250);
   U16264 : OAI22_X1 port map( A1 => n17884, A2 => n16693, B1 => n16784, B2 => 
                           n16694, ZN => n3249);
   U16265 : OAI22_X1 port map( A1 => n17563, A2 => n16691, B1 => n16785, B2 => 
                           n16694, ZN => n3248);
   U16266 : OAI22_X1 port map( A1 => n17564, A2 => n16693, B1 => n16786, B2 => 
                           n16694, ZN => n3247);
   U16267 : OAI22_X1 port map( A1 => n17256, A2 => n16691, B1 => n16787, B2 => 
                           n16694, ZN => n3246);
   U16268 : OAI22_X1 port map( A1 => n17885, A2 => n16691, B1 => n16788, B2 => 
                           n16694, ZN => n3245);
   U16269 : OAI22_X1 port map( A1 => n17565, A2 => n16691, B1 => n16789, B2 => 
                           n16694, ZN => n3244);
   U16270 : OAI22_X1 port map( A1 => n17566, A2 => n16691, B1 => n16790, B2 => 
                           n16694, ZN => n3243);
   U16271 : OAI22_X1 port map( A1 => n17567, A2 => n16691, B1 => n16791, B2 => 
                           n16694, ZN => n3242);
   U16272 : OAI22_X1 port map( A1 => n17257, A2 => n16691, B1 => n16792, B2 => 
                           n16694, ZN => n3241);
   U16273 : OAI22_X1 port map( A1 => n17568, A2 => n16691, B1 => n16793, B2 => 
                           n16694, ZN => n3240);
   U16274 : OAI22_X1 port map( A1 => n18690, A2 => n16693, B1 => n16794, B2 => 
                           n16694, ZN => n3239);
   U16275 : OAI22_X1 port map( A1 => n18925, A2 => n16693, B1 => n16795, B2 => 
                           n16694, ZN => n3238);
   U16276 : OAI22_X1 port map( A1 => n18926, A2 => n16691, B1 => n16796, B2 => 
                           n16694, ZN => n3237);
   U16277 : OAI22_X1 port map( A1 => n18238, A2 => n16691, B1 => n16797, B2 => 
                           n16694, ZN => n3236);
   U16278 : OAI22_X1 port map( A1 => n18927, A2 => n16693, B1 => n16798, B2 => 
                           n16694, ZN => n3235);
   U16279 : OAI22_X1 port map( A1 => n18691, A2 => n16691, B1 => n16799, B2 => 
                           n16694, ZN => n3234);
   U16280 : OAI22_X1 port map( A1 => n18692, A2 => n16693, B1 => n16800, B2 => 
                           n16694, ZN => n3233);
   U16281 : OAI22_X1 port map( A1 => n18693, A2 => n16691, B1 => n16801, B2 => 
                           n16694, ZN => n3232);
   U16282 : OAI22_X1 port map( A1 => n18694, A2 => n16693, B1 => n16802, B2 => 
                           n16694, ZN => n3231);
   U16283 : OAI22_X1 port map( A1 => n18239, A2 => n16693, B1 => n16803, B2 => 
                           n16694, ZN => n3230);
   U16284 : OAI22_X1 port map( A1 => n18928, A2 => n16691, B1 => n16804, B2 => 
                           n16694, ZN => n3229);
   U16285 : OAI22_X1 port map( A1 => n18695, A2 => n16691, B1 => n16805, B2 => 
                           n16692, ZN => n3228);
   U16286 : OAI22_X1 port map( A1 => n18929, A2 => n16693, B1 => n16806, B2 => 
                           n16694, ZN => n3227);
   U16287 : OAI22_X1 port map( A1 => n18696, A2 => n16691, B1 => n16808, B2 => 
                           n16694, ZN => n3226);
   U16288 : OAI22_X1 port map( A1 => n18930, A2 => n16693, B1 => n16810, B2 => 
                           n16692, ZN => n3225);
   U16289 : OAI22_X1 port map( A1 => n18697, A2 => n16691, B1 => n16812, B2 => 
                           n16694, ZN => n3224);
   U16290 : NAND2_X1 port map( A1 => n16734, A2 => n16707, ZN => n16696);
   U16291 : CLKBUF_X2 port map( A => n16696, Z => n16698);
   U16292 : NAND2_X1 port map( A1 => n13731, A2 => n16698, ZN => n16697);
   U16293 : OAI22_X1 port map( A1 => n18011, A2 => n16697, B1 => n16815, B2 => 
                           n16696, ZN => n3223);
   U16294 : CLKBUF_X2 port map( A => n16697, Z => n16695);
   U16295 : OAI22_X1 port map( A1 => n16966, A2 => n16695, B1 => n16816, B2 => 
                           n16698, ZN => n3222);
   U16296 : OAI22_X1 port map( A1 => n16889, A2 => n16697, B1 => n16817, B2 => 
                           n16696, ZN => n3221);
   U16297 : OAI22_X1 port map( A1 => n16967, A2 => n16695, B1 => n16818, B2 => 
                           n16696, ZN => n3220);
   U16298 : OAI22_X1 port map( A1 => n16968, A2 => n16695, B1 => n16819, B2 => 
                           n16698, ZN => n3219);
   U16299 : OAI22_X1 port map( A1 => n16969, A2 => n16695, B1 => n16820, B2 => 
                           n16696, ZN => n3218);
   U16300 : OAI22_X1 port map( A1 => n17108, A2 => n16695, B1 => n16821, B2 => 
                           n16698, ZN => n3217);
   U16301 : OAI22_X1 port map( A1 => n16970, A2 => n16695, B1 => n16822, B2 => 
                           n16698, ZN => n3216);
   U16302 : OAI22_X1 port map( A1 => n16890, A2 => n16695, B1 => n16823, B2 => 
                           n16698, ZN => n3215);
   U16303 : OAI22_X1 port map( A1 => n16891, A2 => n16695, B1 => n16824, B2 => 
                           n16698, ZN => n3214);
   U16304 : OAI22_X1 port map( A1 => n17109, A2 => n16695, B1 => n16825, B2 => 
                           n16698, ZN => n3213);
   U16305 : OAI22_X1 port map( A1 => n16892, A2 => n16695, B1 => n16826, B2 => 
                           n16696, ZN => n3212);
   U16306 : OAI22_X1 port map( A1 => n17569, A2 => n16697, B1 => n16827, B2 => 
                           n16696, ZN => n3211);
   U16307 : OAI22_X1 port map( A1 => n17570, A2 => n16695, B1 => n16828, B2 => 
                           n16698, ZN => n3210);
   U16308 : OAI22_X1 port map( A1 => n17571, A2 => n16695, B1 => n16829, B2 => 
                           n16696, ZN => n3209);
   U16309 : OAI22_X1 port map( A1 => n17572, A2 => n16697, B1 => n16830, B2 => 
                           n16696, ZN => n3208);
   U16310 : OAI22_X1 port map( A1 => n17886, A2 => n16697, B1 => n16831, B2 => 
                           n16696, ZN => n3207);
   U16311 : OAI22_X1 port map( A1 => n17258, A2 => n16695, B1 => n16832, B2 => 
                           n16698, ZN => n3206);
   U16312 : OAI22_X1 port map( A1 => n17259, A2 => n16695, B1 => n16833, B2 => 
                           n16696, ZN => n3205);
   U16313 : OAI22_X1 port map( A1 => n17887, A2 => n16697, B1 => n16834, B2 => 
                           n16696, ZN => n3204);
   U16314 : OAI22_X1 port map( A1 => n17573, A2 => n16697, B1 => n16835, B2 => 
                           n16698, ZN => n3203);
   U16315 : OAI22_X1 port map( A1 => n17574, A2 => n16695, B1 => n16836, B2 => 
                           n16698, ZN => n3202);
   U16316 : OAI22_X1 port map( A1 => n17260, A2 => n16695, B1 => n16837, B2 => 
                           n16698, ZN => n3201);
   U16317 : OAI22_X1 port map( A1 => n17888, A2 => n16695, B1 => n16838, B2 => 
                           n16696, ZN => n3200);
   U16318 : OAI22_X1 port map( A1 => n17575, A2 => n16695, B1 => n16839, B2 => 
                           n16698, ZN => n3199);
   U16319 : OAI22_X1 port map( A1 => n17261, A2 => n16697, B1 => n16840, B2 => 
                           n16696, ZN => n3198);
   U16320 : OAI22_X1 port map( A1 => n17889, A2 => n16695, B1 => n16841, B2 => 
                           n16696, ZN => n3197);
   U16321 : OAI22_X1 port map( A1 => n17262, A2 => n16697, B1 => n16842, B2 => 
                           n16696, ZN => n3196);
   U16322 : OAI22_X1 port map( A1 => n17576, A2 => n16695, B1 => n16843, B2 => 
                           n16696, ZN => n3195);
   U16323 : OAI22_X1 port map( A1 => n17263, A2 => n16697, B1 => n16844, B2 => 
                           n16696, ZN => n3194);
   U16324 : OAI22_X1 port map( A1 => n17890, A2 => n16695, B1 => n16845, B2 => 
                           n16696, ZN => n3193);
   U16325 : OAI22_X1 port map( A1 => n17577, A2 => n16697, B1 => n16846, B2 => 
                           n16696, ZN => n3192);
   U16326 : OAI22_X1 port map( A1 => n17891, A2 => n16695, B1 => n16847, B2 => 
                           n16696, ZN => n3191);
   U16327 : OAI22_X1 port map( A1 => n17892, A2 => n16697, B1 => n16848, B2 => 
                           n16696, ZN => n3190);
   U16328 : OAI22_X1 port map( A1 => n17578, A2 => n16695, B1 => n16849, B2 => 
                           n16696, ZN => n3189);
   U16329 : OAI22_X1 port map( A1 => n17579, A2 => n16697, B1 => n16850, B2 => 
                           n16698, ZN => n3188);
   U16330 : OAI22_X1 port map( A1 => n16893, A2 => n16697, B1 => n16851, B2 => 
                           n16698, ZN => n3187);
   U16331 : OAI22_X1 port map( A1 => n16971, A2 => n16695, B1 => n16852, B2 => 
                           n16698, ZN => n3186);
   U16332 : OAI22_X1 port map( A1 => n16972, A2 => n16697, B1 => n16853, B2 => 
                           n16698, ZN => n3185);
   U16333 : OAI22_X1 port map( A1 => n16973, A2 => n16695, B1 => n16854, B2 => 
                           n16698, ZN => n3184);
   U16334 : OAI22_X1 port map( A1 => n16974, A2 => n16697, B1 => n16855, B2 => 
                           n16698, ZN => n3183);
   U16335 : OAI22_X1 port map( A1 => n16894, A2 => n16695, B1 => n16856, B2 => 
                           n16698, ZN => n3182);
   U16336 : OAI22_X1 port map( A1 => n16975, A2 => n16695, B1 => n16857, B2 => 
                           n16698, ZN => n3181);
   U16337 : OAI22_X1 port map( A1 => n16976, A2 => n16695, B1 => n16858, B2 => 
                           n16698, ZN => n3180);
   U16338 : OAI22_X1 port map( A1 => n16977, A2 => n16695, B1 => n16859, B2 => 
                           n16698, ZN => n3179);
   U16339 : OAI22_X1 port map( A1 => n17110, A2 => n16695, B1 => n16860, B2 => 
                           n16698, ZN => n3178);
   U16340 : OAI22_X1 port map( A1 => n17111, A2 => n16695, B1 => n16861, B2 => 
                           n16698, ZN => n3177);
   U16341 : OAI22_X1 port map( A1 => n16978, A2 => n16695, B1 => n16862, B2 => 
                           n16698, ZN => n3176);
   U16342 : OAI22_X1 port map( A1 => n17893, A2 => n16697, B1 => n16863, B2 => 
                           n16698, ZN => n3175);
   U16343 : OAI22_X1 port map( A1 => n17894, A2 => n16697, B1 => n16864, B2 => 
                           n16698, ZN => n3174);
   U16344 : OAI22_X1 port map( A1 => n17580, A2 => n16695, B1 => n16865, B2 => 
                           n16698, ZN => n3173);
   U16345 : OAI22_X1 port map( A1 => n17581, A2 => n16695, B1 => n16866, B2 => 
                           n16698, ZN => n3172);
   U16346 : OAI22_X1 port map( A1 => n17895, A2 => n16697, B1 => n16867, B2 => 
                           n16698, ZN => n3171);
   U16347 : OAI22_X1 port map( A1 => n17264, A2 => n16695, B1 => n16868, B2 => 
                           n16698, ZN => n3170);
   U16348 : OAI22_X1 port map( A1 => n17582, A2 => n16697, B1 => n16869, B2 => 
                           n16698, ZN => n3169);
   U16349 : OAI22_X1 port map( A1 => n17265, A2 => n16695, B1 => n16870, B2 => 
                           n16698, ZN => n3168);
   U16350 : OAI22_X1 port map( A1 => n17896, A2 => n16697, B1 => n16871, B2 => 
                           n16698, ZN => n3167);
   U16351 : OAI22_X1 port map( A1 => n17897, A2 => n16697, B1 => n16872, B2 => 
                           n16698, ZN => n3166);
   U16352 : OAI22_X1 port map( A1 => n17583, A2 => n16695, B1 => n16873, B2 => 
                           n16698, ZN => n3165);
   U16353 : OAI22_X1 port map( A1 => n17584, A2 => n16695, B1 => n16874, B2 => 
                           n16696, ZN => n3164);
   U16354 : OAI22_X1 port map( A1 => n17585, A2 => n16697, B1 => n16875, B2 => 
                           n16698, ZN => n3163);
   U16355 : OAI22_X1 port map( A1 => n17898, A2 => n16695, B1 => n16876, B2 => 
                           n16698, ZN => n3162);
   U16356 : OAI22_X1 port map( A1 => n17899, A2 => n16697, B1 => n16878, B2 => 
                           n16696, ZN => n3161);
   U16357 : OAI22_X1 port map( A1 => n17900, A2 => n16695, B1 => n16881, B2 => 
                           n16698, ZN => n3160);
   U16358 : NAND2_X1 port map( A1 => n16739, A2 => n16707, ZN => n16700);
   U16359 : CLKBUF_X2 port map( A => n16700, Z => n16702);
   U16360 : NAND2_X1 port map( A1 => n13731, A2 => n16702, ZN => n16701);
   U16361 : OAI22_X1 port map( A1 => n18012, A2 => n16701, B1 => n16745, B2 => 
                           n16700, ZN => n3159);
   U16362 : CLKBUF_X2 port map( A => n16701, Z => n16699);
   U16363 : OAI22_X1 port map( A1 => n16895, A2 => n16699, B1 => n16816, B2 => 
                           n16702, ZN => n3158);
   U16364 : OAI22_X1 port map( A1 => n16979, A2 => n16701, B1 => n16817, B2 => 
                           n16700, ZN => n3157);
   U16365 : OAI22_X1 port map( A1 => n16896, A2 => n16699, B1 => n16818, B2 => 
                           n16700, ZN => n3156);
   U16366 : OAI22_X1 port map( A1 => n16980, A2 => n16699, B1 => n16819, B2 => 
                           n16702, ZN => n3155);
   U16367 : OAI22_X1 port map( A1 => n16981, A2 => n16699, B1 => n16820, B2 => 
                           n16700, ZN => n3154);
   U16368 : OAI22_X1 port map( A1 => n16982, A2 => n16699, B1 => n16821, B2 => 
                           n16702, ZN => n3153);
   U16369 : OAI22_X1 port map( A1 => n16983, A2 => n16699, B1 => n16822, B2 => 
                           n16702, ZN => n3152);
   U16370 : OAI22_X1 port map( A1 => n16984, A2 => n16699, B1 => n16823, B2 => 
                           n16702, ZN => n3151);
   U16371 : OAI22_X1 port map( A1 => n16897, A2 => n16699, B1 => n16824, B2 => 
                           n16702, ZN => n3150);
   U16372 : OAI22_X1 port map( A1 => n16985, A2 => n16699, B1 => n16825, B2 => 
                           n16702, ZN => n3149);
   U16373 : OAI22_X1 port map( A1 => n16898, A2 => n16699, B1 => n16826, B2 => 
                           n16700, ZN => n3148);
   U16374 : OAI22_X1 port map( A1 => n17586, A2 => n16701, B1 => n16827, B2 => 
                           n16700, ZN => n3147);
   U16375 : OAI22_X1 port map( A1 => n17266, A2 => n16699, B1 => n16828, B2 => 
                           n16702, ZN => n3146);
   U16376 : OAI22_X1 port map( A1 => n17587, A2 => n16699, B1 => n16829, B2 => 
                           n16700, ZN => n3145);
   U16377 : OAI22_X1 port map( A1 => n17267, A2 => n16701, B1 => n16830, B2 => 
                           n16700, ZN => n3144);
   U16378 : OAI22_X1 port map( A1 => n17588, A2 => n16701, B1 => n16831, B2 => 
                           n16700, ZN => n3143);
   U16379 : OAI22_X1 port map( A1 => n17589, A2 => n16699, B1 => n16832, B2 => 
                           n16702, ZN => n3142);
   U16380 : OAI22_X1 port map( A1 => n17590, A2 => n16699, B1 => n16833, B2 => 
                           n16700, ZN => n3141);
   U16381 : OAI22_X1 port map( A1 => n17591, A2 => n16701, B1 => n16834, B2 => 
                           n16700, ZN => n3140);
   U16382 : OAI22_X1 port map( A1 => n17268, A2 => n16701, B1 => n16835, B2 => 
                           n16702, ZN => n3139);
   U16383 : OAI22_X1 port map( A1 => n17592, A2 => n16699, B1 => n16836, B2 => 
                           n16702, ZN => n3138);
   U16384 : OAI22_X1 port map( A1 => n17269, A2 => n16699, B1 => n16837, B2 => 
                           n16702, ZN => n3137);
   U16385 : OAI22_X1 port map( A1 => n17593, A2 => n16699, B1 => n16838, B2 => 
                           n16700, ZN => n3136);
   U16386 : OAI22_X1 port map( A1 => n17594, A2 => n16699, B1 => n16839, B2 => 
                           n16702, ZN => n3135);
   U16387 : OAI22_X1 port map( A1 => n17270, A2 => n16701, B1 => n16840, B2 => 
                           n16700, ZN => n3134);
   U16388 : OAI22_X1 port map( A1 => n17271, A2 => n16699, B1 => n16841, B2 => 
                           n16700, ZN => n3133);
   U16389 : OAI22_X1 port map( A1 => n17272, A2 => n16701, B1 => n16842, B2 => 
                           n16700, ZN => n3132);
   U16390 : OAI22_X1 port map( A1 => n17595, A2 => n16699, B1 => n16843, B2 => 
                           n16700, ZN => n3131);
   U16391 : OAI22_X1 port map( A1 => n17596, A2 => n16701, B1 => n16844, B2 => 
                           n16700, ZN => n3130);
   U16392 : OAI22_X1 port map( A1 => n17597, A2 => n16699, B1 => n16845, B2 => 
                           n16700, ZN => n3129);
   U16393 : OAI22_X1 port map( A1 => n17598, A2 => n16701, B1 => n16846, B2 => 
                           n16700, ZN => n3128);
   U16394 : OAI22_X1 port map( A1 => n17273, A2 => n16699, B1 => n16847, B2 => 
                           n16700, ZN => n3127);
   U16395 : OAI22_X1 port map( A1 => n17274, A2 => n16701, B1 => n16848, B2 => 
                           n16700, ZN => n3126);
   U16396 : OAI22_X1 port map( A1 => n17275, A2 => n16699, B1 => n16849, B2 => 
                           n16700, ZN => n3125);
   U16397 : OAI22_X1 port map( A1 => n17276, A2 => n16701, B1 => n16850, B2 => 
                           n16702, ZN => n3124);
   U16398 : OAI22_X1 port map( A1 => n16986, A2 => n16701, B1 => n16851, B2 => 
                           n16702, ZN => n3123);
   U16399 : OAI22_X1 port map( A1 => n16899, A2 => n16699, B1 => n16852, B2 => 
                           n16702, ZN => n3122);
   U16400 : OAI22_X1 port map( A1 => n16987, A2 => n16701, B1 => n16853, B2 => 
                           n16702, ZN => n3121);
   U16401 : OAI22_X1 port map( A1 => n16900, A2 => n16699, B1 => n16854, B2 => 
                           n16702, ZN => n3120);
   U16402 : OAI22_X1 port map( A1 => n16901, A2 => n16701, B1 => n16855, B2 => 
                           n16702, ZN => n3119);
   U16403 : OAI22_X1 port map( A1 => n16902, A2 => n16699, B1 => n16856, B2 => 
                           n16702, ZN => n3118);
   U16404 : OAI22_X1 port map( A1 => n16988, A2 => n16699, B1 => n16857, B2 => 
                           n16702, ZN => n3117);
   U16405 : OAI22_X1 port map( A1 => n16903, A2 => n16699, B1 => n16858, B2 => 
                           n16702, ZN => n3116);
   U16406 : OAI22_X1 port map( A1 => n16989, A2 => n16699, B1 => n16859, B2 => 
                           n16702, ZN => n3115);
   U16407 : OAI22_X1 port map( A1 => n16990, A2 => n16699, B1 => n16860, B2 => 
                           n16702, ZN => n3114);
   U16408 : OAI22_X1 port map( A1 => n16991, A2 => n16699, B1 => n16861, B2 => 
                           n16702, ZN => n3113);
   U16409 : OAI22_X1 port map( A1 => n16904, A2 => n16699, B1 => n16862, B2 => 
                           n16702, ZN => n3112);
   U16410 : OAI22_X1 port map( A1 => n17599, A2 => n16701, B1 => n16863, B2 => 
                           n16702, ZN => n3111);
   U16411 : OAI22_X1 port map( A1 => n17600, A2 => n16701, B1 => n16864, B2 => 
                           n16702, ZN => n3110);
   U16412 : OAI22_X1 port map( A1 => n17601, A2 => n16699, B1 => n16865, B2 => 
                           n16702, ZN => n3109);
   U16413 : OAI22_X1 port map( A1 => n17602, A2 => n16699, B1 => n16866, B2 => 
                           n16702, ZN => n3108);
   U16414 : OAI22_X1 port map( A1 => n17603, A2 => n16701, B1 => n16867, B2 => 
                           n16702, ZN => n3107);
   U16415 : OAI22_X1 port map( A1 => n17604, A2 => n16699, B1 => n16868, B2 => 
                           n16702, ZN => n3106);
   U16416 : OAI22_X1 port map( A1 => n17605, A2 => n16701, B1 => n16869, B2 => 
                           n16702, ZN => n3105);
   U16417 : OAI22_X1 port map( A1 => n17277, A2 => n16699, B1 => n16870, B2 => 
                           n16702, ZN => n3104);
   U16418 : OAI22_X1 port map( A1 => n17606, A2 => n16701, B1 => n16871, B2 => 
                           n16702, ZN => n3103);
   U16419 : OAI22_X1 port map( A1 => n17607, A2 => n16701, B1 => n16872, B2 => 
                           n16702, ZN => n3102);
   U16420 : OAI22_X1 port map( A1 => n17608, A2 => n16699, B1 => n16873, B2 => 
                           n16702, ZN => n3101);
   U16421 : OAI22_X1 port map( A1 => n17278, A2 => n16699, B1 => n16874, B2 => 
                           n16700, ZN => n3100);
   U16422 : OAI22_X1 port map( A1 => n17279, A2 => n16701, B1 => n16875, B2 => 
                           n16702, ZN => n3099);
   U16423 : OAI22_X1 port map( A1 => n17609, A2 => n16699, B1 => n16876, B2 => 
                           n16702, ZN => n3098);
   U16424 : OAI22_X1 port map( A1 => n17610, A2 => n16701, B1 => n16878, B2 => 
                           n16700, ZN => n3097);
   U16425 : OAI22_X1 port map( A1 => n17611, A2 => n16699, B1 => n16881, B2 => 
                           n16702, ZN => n3096);
   U16426 : NAND2_X1 port map( A1 => n16744, A2 => n16707, ZN => n16704);
   U16427 : CLKBUF_X2 port map( A => n16704, Z => n16706);
   U16428 : NAND2_X1 port map( A1 => n13731, A2 => n16706, ZN => n16705);
   U16429 : OAI22_X1 port map( A1 => n18240, A2 => n16705, B1 => n16815, B2 => 
                           n16704, ZN => n3095);
   U16430 : CLKBUF_X2 port map( A => n16705, Z => n16703);
   U16431 : OAI22_X1 port map( A1 => n16905, A2 => n16703, B1 => n16746, B2 => 
                           n16706, ZN => n3094);
   U16432 : OAI22_X1 port map( A1 => n16906, A2 => n16705, B1 => n16747, B2 => 
                           n16704, ZN => n3093);
   U16433 : OAI22_X1 port map( A1 => n16992, A2 => n16703, B1 => n16748, B2 => 
                           n16704, ZN => n3092);
   U16434 : OAI22_X1 port map( A1 => n16993, A2 => n16703, B1 => n16749, B2 => 
                           n16706, ZN => n3091);
   U16435 : OAI22_X1 port map( A1 => n16994, A2 => n16703, B1 => n16750, B2 => 
                           n16704, ZN => n3090);
   U16436 : OAI22_X1 port map( A1 => n16995, A2 => n16703, B1 => n16751, B2 => 
                           n16706, ZN => n3089);
   U16437 : OAI22_X1 port map( A1 => n16996, A2 => n16703, B1 => n16752, B2 => 
                           n16706, ZN => n3088);
   U16438 : OAI22_X1 port map( A1 => n16997, A2 => n16703, B1 => n16753, B2 => 
                           n16706, ZN => n3087);
   U16439 : OAI22_X1 port map( A1 => n16907, A2 => n16703, B1 => n16754, B2 => 
                           n16706, ZN => n3086);
   U16440 : OAI22_X1 port map( A1 => n17112, A2 => n16703, B1 => n16755, B2 => 
                           n16706, ZN => n3085);
   U16441 : OAI22_X1 port map( A1 => n16998, A2 => n16703, B1 => n16756, B2 => 
                           n16704, ZN => n3084);
   U16442 : OAI22_X1 port map( A1 => n17280, A2 => n16705, B1 => n16757, B2 => 
                           n16704, ZN => n3083);
   U16443 : OAI22_X1 port map( A1 => n17281, A2 => n16703, B1 => n16758, B2 => 
                           n16706, ZN => n3082);
   U16444 : OAI22_X1 port map( A1 => n17282, A2 => n16703, B1 => n16759, B2 => 
                           n16704, ZN => n3081);
   U16445 : OAI22_X1 port map( A1 => n17283, A2 => n16705, B1 => n16760, B2 => 
                           n16704, ZN => n3080);
   U16446 : OAI22_X1 port map( A1 => n17612, A2 => n16705, B1 => n16761, B2 => 
                           n16704, ZN => n3079);
   U16447 : OAI22_X1 port map( A1 => n17284, A2 => n16703, B1 => n16762, B2 => 
                           n16706, ZN => n3078);
   U16448 : OAI22_X1 port map( A1 => n17613, A2 => n16703, B1 => n16763, B2 => 
                           n16704, ZN => n3077);
   U16449 : OAI22_X1 port map( A1 => n17285, A2 => n16705, B1 => n16764, B2 => 
                           n16704, ZN => n3076);
   U16450 : OAI22_X1 port map( A1 => n17286, A2 => n16705, B1 => n16765, B2 => 
                           n16706, ZN => n3075);
   U16451 : OAI22_X1 port map( A1 => n17614, A2 => n16703, B1 => n16766, B2 => 
                           n16706, ZN => n3074);
   U16452 : OAI22_X1 port map( A1 => n17615, A2 => n16703, B1 => n16767, B2 => 
                           n16706, ZN => n3073);
   U16453 : OAI22_X1 port map( A1 => n17616, A2 => n16703, B1 => n16768, B2 => 
                           n16704, ZN => n3072);
   U16454 : OAI22_X1 port map( A1 => n17287, A2 => n16703, B1 => n16769, B2 => 
                           n16706, ZN => n3071);
   U16455 : OAI22_X1 port map( A1 => n17288, A2 => n16705, B1 => n16770, B2 => 
                           n16704, ZN => n3070);
   U16456 : OAI22_X1 port map( A1 => n17289, A2 => n16703, B1 => n16771, B2 => 
                           n16704, ZN => n3069);
   U16457 : OAI22_X1 port map( A1 => n17617, A2 => n16705, B1 => n16772, B2 => 
                           n16704, ZN => n3068);
   U16458 : OAI22_X1 port map( A1 => n17618, A2 => n16703, B1 => n16773, B2 => 
                           n16704, ZN => n3067);
   U16459 : OAI22_X1 port map( A1 => n17290, A2 => n16705, B1 => n16774, B2 => 
                           n16704, ZN => n3066);
   U16460 : OAI22_X1 port map( A1 => n17291, A2 => n16703, B1 => n16775, B2 => 
                           n16704, ZN => n3065);
   U16461 : OAI22_X1 port map( A1 => n17619, A2 => n16705, B1 => n16776, B2 => 
                           n16704, ZN => n3064);
   U16462 : OAI22_X1 port map( A1 => n17620, A2 => n16703, B1 => n16777, B2 => 
                           n16704, ZN => n3063);
   U16463 : OAI22_X1 port map( A1 => n17621, A2 => n16705, B1 => n16778, B2 => 
                           n16704, ZN => n3062);
   U16464 : OAI22_X1 port map( A1 => n17292, A2 => n16703, B1 => n16779, B2 => 
                           n16704, ZN => n3061);
   U16465 : OAI22_X1 port map( A1 => n17622, A2 => n16705, B1 => n16781, B2 => 
                           n16706, ZN => n3060);
   U16466 : OAI22_X1 port map( A1 => n16908, A2 => n16705, B1 => n16782, B2 => 
                           n16706, ZN => n3059);
   U16467 : OAI22_X1 port map( A1 => n16909, A2 => n16703, B1 => n16783, B2 => 
                           n16706, ZN => n3058);
   U16468 : OAI22_X1 port map( A1 => n16999, A2 => n16705, B1 => n16784, B2 => 
                           n16706, ZN => n3057);
   U16469 : OAI22_X1 port map( A1 => n17000, A2 => n16703, B1 => n16785, B2 => 
                           n16706, ZN => n3056);
   U16470 : OAI22_X1 port map( A1 => n16910, A2 => n16705, B1 => n16786, B2 => 
                           n16706, ZN => n3055);
   U16471 : OAI22_X1 port map( A1 => n17001, A2 => n16703, B1 => n16787, B2 => 
                           n16706, ZN => n3054);
   U16472 : OAI22_X1 port map( A1 => n16911, A2 => n16703, B1 => n16788, B2 => 
                           n16706, ZN => n3053);
   U16473 : OAI22_X1 port map( A1 => n16912, A2 => n16703, B1 => n16789, B2 => 
                           n16706, ZN => n3052);
   U16474 : OAI22_X1 port map( A1 => n17113, A2 => n16703, B1 => n16790, B2 => 
                           n16706, ZN => n3051);
   U16475 : OAI22_X1 port map( A1 => n16913, A2 => n16703, B1 => n16791, B2 => 
                           n16706, ZN => n3050);
   U16476 : OAI22_X1 port map( A1 => n16914, A2 => n16703, B1 => n16792, B2 => 
                           n16706, ZN => n3049);
   U16477 : OAI22_X1 port map( A1 => n17002, A2 => n16703, B1 => n16793, B2 => 
                           n16706, ZN => n3048);
   U16478 : OAI22_X1 port map( A1 => n17623, A2 => n16705, B1 => n16794, B2 => 
                           n16706, ZN => n3047);
   U16479 : OAI22_X1 port map( A1 => n17293, A2 => n16705, B1 => n16795, B2 => 
                           n16706, ZN => n3046);
   U16480 : OAI22_X1 port map( A1 => n17624, A2 => n16703, B1 => n16796, B2 => 
                           n16706, ZN => n3045);
   U16481 : OAI22_X1 port map( A1 => n17294, A2 => n16703, B1 => n16797, B2 => 
                           n16706, ZN => n3044);
   U16482 : OAI22_X1 port map( A1 => n17295, A2 => n16705, B1 => n16798, B2 => 
                           n16706, ZN => n3043);
   U16483 : OAI22_X1 port map( A1 => n17625, A2 => n16703, B1 => n16799, B2 => 
                           n16706, ZN => n3042);
   U16484 : OAI22_X1 port map( A1 => n17296, A2 => n16705, B1 => n16800, B2 => 
                           n16706, ZN => n3041);
   U16485 : OAI22_X1 port map( A1 => n17297, A2 => n16703, B1 => n16801, B2 => 
                           n16706, ZN => n3040);
   U16486 : OAI22_X1 port map( A1 => n17626, A2 => n16705, B1 => n16802, B2 => 
                           n16706, ZN => n3039);
   U16487 : OAI22_X1 port map( A1 => n17298, A2 => n16705, B1 => n16803, B2 => 
                           n16706, ZN => n3038);
   U16488 : OAI22_X1 port map( A1 => n17627, A2 => n16703, B1 => n16804, B2 => 
                           n16706, ZN => n3037);
   U16489 : OAI22_X1 port map( A1 => n17299, A2 => n16703, B1 => n16805, B2 => 
                           n16704, ZN => n3036);
   U16490 : OAI22_X1 port map( A1 => n17628, A2 => n16705, B1 => n16806, B2 => 
                           n16706, ZN => n3035);
   U16491 : OAI22_X1 port map( A1 => n17300, A2 => n16703, B1 => n16808, B2 => 
                           n16706, ZN => n3034);
   U16492 : OAI22_X1 port map( A1 => n17301, A2 => n16705, B1 => n16810, B2 => 
                           n16704, ZN => n3033);
   U16493 : OAI22_X1 port map( A1 => n17629, A2 => n16703, B1 => n16812, B2 => 
                           n16706, ZN => n3032);
   U16494 : NAND2_X1 port map( A1 => n16814, A2 => n16707, ZN => n16709);
   U16495 : CLKBUF_X2 port map( A => n16709, Z => n16711);
   U16496 : NAND2_X1 port map( A1 => n13731, A2 => n16711, ZN => n16710);
   U16497 : OAI22_X1 port map( A1 => n18698, A2 => n16710, B1 => n16815, B2 => 
                           n16709, ZN => n3031);
   U16498 : CLKBUF_X2 port map( A => n16710, Z => n16708);
   U16499 : OAI22_X1 port map( A1 => n17003, A2 => n16708, B1 => n16816, B2 => 
                           n16711, ZN => n3030);
   U16500 : OAI22_X1 port map( A1 => n17114, A2 => n16710, B1 => n16817, B2 => 
                           n16709, ZN => n3029);
   U16501 : OAI22_X1 port map( A1 => n17004, A2 => n16708, B1 => n16818, B2 => 
                           n16709, ZN => n3028);
   U16502 : OAI22_X1 port map( A1 => n17005, A2 => n16708, B1 => n16819, B2 => 
                           n16711, ZN => n3027);
   U16503 : OAI22_X1 port map( A1 => n17006, A2 => n16708, B1 => n16820, B2 => 
                           n16709, ZN => n3026);
   U16504 : OAI22_X1 port map( A1 => n17115, A2 => n16708, B1 => n16821, B2 => 
                           n16711, ZN => n3025);
   U16505 : OAI22_X1 port map( A1 => n17007, A2 => n16708, B1 => n16822, B2 => 
                           n16711, ZN => n3024);
   U16506 : OAI22_X1 port map( A1 => n16915, A2 => n16708, B1 => n16823, B2 => 
                           n16711, ZN => n3023);
   U16507 : OAI22_X1 port map( A1 => n17008, A2 => n16708, B1 => n16824, B2 => 
                           n16711, ZN => n3022);
   U16508 : OAI22_X1 port map( A1 => n17009, A2 => n16708, B1 => n16825, B2 => 
                           n16711, ZN => n3021);
   U16509 : OAI22_X1 port map( A1 => n17116, A2 => n16708, B1 => n16826, B2 => 
                           n16709, ZN => n3020);
   U16510 : OAI22_X1 port map( A1 => n17630, A2 => n16710, B1 => n16827, B2 => 
                           n16709, ZN => n3019);
   U16511 : OAI22_X1 port map( A1 => n17631, A2 => n16708, B1 => n16828, B2 => 
                           n16711, ZN => n3018);
   U16512 : OAI22_X1 port map( A1 => n17632, A2 => n16708, B1 => n16829, B2 => 
                           n16709, ZN => n3017);
   U16513 : OAI22_X1 port map( A1 => n17633, A2 => n16710, B1 => n16830, B2 => 
                           n16709, ZN => n3016);
   U16514 : OAI22_X1 port map( A1 => n17901, A2 => n16710, B1 => n16831, B2 => 
                           n16709, ZN => n3015);
   U16515 : OAI22_X1 port map( A1 => n17902, A2 => n16708, B1 => n16832, B2 => 
                           n16711, ZN => n3014);
   U16516 : OAI22_X1 port map( A1 => n17302, A2 => n16708, B1 => n16833, B2 => 
                           n16709, ZN => n3013);
   U16517 : OAI22_X1 port map( A1 => n17634, A2 => n16710, B1 => n16834, B2 => 
                           n16709, ZN => n3012);
   U16518 : OAI22_X1 port map( A1 => n17635, A2 => n16710, B1 => n16835, B2 => 
                           n16711, ZN => n3011);
   U16519 : OAI22_X1 port map( A1 => n17903, A2 => n16708, B1 => n16836, B2 => 
                           n16711, ZN => n3010);
   U16520 : OAI22_X1 port map( A1 => n17904, A2 => n16708, B1 => n16837, B2 => 
                           n16711, ZN => n3009);
   U16521 : OAI22_X1 port map( A1 => n17303, A2 => n16708, B1 => n16838, B2 => 
                           n16709, ZN => n3008);
   U16522 : OAI22_X1 port map( A1 => n17636, A2 => n16708, B1 => n16839, B2 => 
                           n16711, ZN => n3007);
   U16523 : OAI22_X1 port map( A1 => n17637, A2 => n16710, B1 => n16840, B2 => 
                           n16709, ZN => n3006);
   U16524 : OAI22_X1 port map( A1 => n17905, A2 => n16708, B1 => n16841, B2 => 
                           n16709, ZN => n3005);
   U16525 : OAI22_X1 port map( A1 => n17906, A2 => n16710, B1 => n16842, B2 => 
                           n16709, ZN => n3004);
   U16526 : OAI22_X1 port map( A1 => n17907, A2 => n16708, B1 => n16843, B2 => 
                           n16709, ZN => n3003);
   U16527 : OAI22_X1 port map( A1 => n17304, A2 => n16710, B1 => n16844, B2 => 
                           n16709, ZN => n3002);
   U16528 : OAI22_X1 port map( A1 => n17638, A2 => n16708, B1 => n16845, B2 => 
                           n16709, ZN => n3001);
   U16529 : OAI22_X1 port map( A1 => n17305, A2 => n16710, B1 => n16846, B2 => 
                           n16709, ZN => n3000);
   U16530 : OAI22_X1 port map( A1 => n17908, A2 => n16708, B1 => n16847, B2 => 
                           n16709, ZN => n2999);
   U16531 : OAI22_X1 port map( A1 => n17909, A2 => n16710, B1 => n16848, B2 => 
                           n16709, ZN => n2998);
   U16532 : OAI22_X1 port map( A1 => n17306, A2 => n16708, B1 => n16849, B2 => 
                           n16709, ZN => n2997);
   U16533 : OAI22_X1 port map( A1 => n17639, A2 => n16710, B1 => n16850, B2 => 
                           n16711, ZN => n2996);
   U16534 : OAI22_X1 port map( A1 => n17010, A2 => n16710, B1 => n16851, B2 => 
                           n16711, ZN => n2995);
   U16535 : OAI22_X1 port map( A1 => n17011, A2 => n16708, B1 => n16852, B2 => 
                           n16711, ZN => n2994);
   U16536 : OAI22_X1 port map( A1 => n16916, A2 => n16710, B1 => n16853, B2 => 
                           n16711, ZN => n2993);
   U16537 : OAI22_X1 port map( A1 => n16917, A2 => n16708, B1 => n16854, B2 => 
                           n16711, ZN => n2992);
   U16538 : OAI22_X1 port map( A1 => n16918, A2 => n16710, B1 => n16855, B2 => 
                           n16711, ZN => n2991);
   U16539 : OAI22_X1 port map( A1 => n17117, A2 => n16708, B1 => n16856, B2 => 
                           n16711, ZN => n2990);
   U16540 : OAI22_X1 port map( A1 => n17012, A2 => n16708, B1 => n16857, B2 => 
                           n16711, ZN => n2989);
   U16541 : OAI22_X1 port map( A1 => n17118, A2 => n16708, B1 => n16858, B2 => 
                           n16711, ZN => n2988);
   U16542 : OAI22_X1 port map( A1 => n17119, A2 => n16708, B1 => n16859, B2 => 
                           n16711, ZN => n2987);
   U16543 : OAI22_X1 port map( A1 => n17013, A2 => n16708, B1 => n16860, B2 => 
                           n16711, ZN => n2986);
   U16544 : OAI22_X1 port map( A1 => n17120, A2 => n16708, B1 => n16861, B2 => 
                           n16711, ZN => n2985);
   U16545 : OAI22_X1 port map( A1 => n17014, A2 => n16708, B1 => n16862, B2 => 
                           n16711, ZN => n2984);
   U16546 : OAI22_X1 port map( A1 => n17640, A2 => n16710, B1 => n16863, B2 => 
                           n16711, ZN => n2983);
   U16547 : OAI22_X1 port map( A1 => n17641, A2 => n16710, B1 => n16864, B2 => 
                           n16711, ZN => n2982);
   U16548 : OAI22_X1 port map( A1 => n17910, A2 => n16708, B1 => n16865, B2 => 
                           n16711, ZN => n2981);
   U16549 : OAI22_X1 port map( A1 => n17642, A2 => n16708, B1 => n16866, B2 => 
                           n16711, ZN => n2980);
   U16550 : OAI22_X1 port map( A1 => n17643, A2 => n16710, B1 => n16867, B2 => 
                           n16711, ZN => n2979);
   U16551 : OAI22_X1 port map( A1 => n17644, A2 => n16708, B1 => n16868, B2 => 
                           n16711, ZN => n2978);
   U16552 : OAI22_X1 port map( A1 => n17645, A2 => n16710, B1 => n16869, B2 => 
                           n16711, ZN => n2977);
   U16553 : OAI22_X1 port map( A1 => n17307, A2 => n16708, B1 => n16870, B2 => 
                           n16711, ZN => n2976);
   U16554 : OAI22_X1 port map( A1 => n17646, A2 => n16710, B1 => n16871, B2 => 
                           n16711, ZN => n2975);
   U16555 : OAI22_X1 port map( A1 => n17911, A2 => n16710, B1 => n16872, B2 => 
                           n16711, ZN => n2974);
   U16556 : OAI22_X1 port map( A1 => n17308, A2 => n16708, B1 => n16873, B2 => 
                           n16711, ZN => n2973);
   U16557 : OAI22_X1 port map( A1 => n17647, A2 => n16708, B1 => n16874, B2 => 
                           n16709, ZN => n2972);
   U16558 : OAI22_X1 port map( A1 => n17309, A2 => n16710, B1 => n16875, B2 => 
                           n16711, ZN => n2971);
   U16559 : OAI22_X1 port map( A1 => n17310, A2 => n16708, B1 => n16876, B2 => 
                           n16711, ZN => n2970);
   U16560 : OAI22_X1 port map( A1 => n17648, A2 => n16710, B1 => n16878, B2 => 
                           n16709, ZN => n2969);
   U16561 : OAI22_X1 port map( A1 => n17649, A2 => n16708, B1 => n16881, B2 => 
                           n16711, ZN => n2968);
   U16562 : NOR2_X1 port map( A1 => n16713, A2 => n16712, ZN => n16813);
   U16563 : NAND2_X1 port map( A1 => n16714, A2 => n16813, ZN => n16716);
   U16564 : CLKBUF_X2 port map( A => n16716, Z => n16718);
   U16565 : NAND2_X1 port map( A1 => n13731, A2 => n16718, ZN => n16717);
   U16566 : OAI22_X1 port map( A1 => n18013, A2 => n16717, B1 => n16745, B2 => 
                           n16716, ZN => n2967);
   U16567 : CLKBUF_X2 port map( A => n16717, Z => n16715);
   U16568 : OAI22_X1 port map( A1 => n17015, A2 => n16715, B1 => n16746, B2 => 
                           n16718, ZN => n2966);
   U16569 : OAI22_X1 port map( A1 => n17121, A2 => n16717, B1 => n16747, B2 => 
                           n16716, ZN => n2965);
   U16570 : OAI22_X1 port map( A1 => n17122, A2 => n16715, B1 => n16748, B2 => 
                           n16716, ZN => n2964);
   U16571 : OAI22_X1 port map( A1 => n17123, A2 => n16715, B1 => n16749, B2 => 
                           n16718, ZN => n2963);
   U16572 : OAI22_X1 port map( A1 => n16919, A2 => n16715, B1 => n16750, B2 => 
                           n16716, ZN => n2962);
   U16573 : OAI22_X1 port map( A1 => n17016, A2 => n16715, B1 => n16751, B2 => 
                           n16718, ZN => n2961);
   U16574 : OAI22_X1 port map( A1 => n16920, A2 => n16715, B1 => n16752, B2 => 
                           n16718, ZN => n2960);
   U16575 : OAI22_X1 port map( A1 => n17124, A2 => n16715, B1 => n16753, B2 => 
                           n16718, ZN => n2959);
   U16576 : OAI22_X1 port map( A1 => n17125, A2 => n16715, B1 => n16754, B2 => 
                           n16718, ZN => n2958);
   U16577 : OAI22_X1 port map( A1 => n16921, A2 => n16715, B1 => n16755, B2 => 
                           n16718, ZN => n2957);
   U16578 : OAI22_X1 port map( A1 => n17017, A2 => n16715, B1 => n16756, B2 => 
                           n16716, ZN => n2956);
   U16579 : OAI22_X1 port map( A1 => n17650, A2 => n16717, B1 => n16757, B2 => 
                           n16716, ZN => n2955);
   U16580 : OAI22_X1 port map( A1 => n17651, A2 => n16715, B1 => n16758, B2 => 
                           n16718, ZN => n2954);
   U16581 : OAI22_X1 port map( A1 => n17912, A2 => n16715, B1 => n16759, B2 => 
                           n16716, ZN => n2953);
   U16582 : OAI22_X1 port map( A1 => n17652, A2 => n16717, B1 => n16760, B2 => 
                           n16716, ZN => n2952);
   U16583 : OAI22_X1 port map( A1 => n17311, A2 => n16717, B1 => n16761, B2 => 
                           n16716, ZN => n2951);
   U16584 : OAI22_X1 port map( A1 => n17653, A2 => n16715, B1 => n16762, B2 => 
                           n16718, ZN => n2950);
   U16585 : OAI22_X1 port map( A1 => n17654, A2 => n16715, B1 => n16763, B2 => 
                           n16716, ZN => n2949);
   U16586 : OAI22_X1 port map( A1 => n17312, A2 => n16717, B1 => n16764, B2 => 
                           n16716, ZN => n2948);
   U16587 : OAI22_X1 port map( A1 => n17913, A2 => n16717, B1 => n16765, B2 => 
                           n16718, ZN => n2947);
   U16588 : OAI22_X1 port map( A1 => n17313, A2 => n16715, B1 => n16766, B2 => 
                           n16718, ZN => n2946);
   U16589 : OAI22_X1 port map( A1 => n17314, A2 => n16715, B1 => n16767, B2 => 
                           n16718, ZN => n2945);
   U16590 : OAI22_X1 port map( A1 => n17655, A2 => n16715, B1 => n16768, B2 => 
                           n16716, ZN => n2944);
   U16591 : OAI22_X1 port map( A1 => n17656, A2 => n16715, B1 => n16769, B2 => 
                           n16718, ZN => n2943);
   U16592 : OAI22_X1 port map( A1 => n17914, A2 => n16717, B1 => n16770, B2 => 
                           n16716, ZN => n2942);
   U16593 : OAI22_X1 port map( A1 => n17315, A2 => n16715, B1 => n16771, B2 => 
                           n16716, ZN => n2941);
   U16594 : OAI22_X1 port map( A1 => n17316, A2 => n16717, B1 => n16772, B2 => 
                           n16716, ZN => n2940);
   U16595 : OAI22_X1 port map( A1 => n17657, A2 => n16715, B1 => n16773, B2 => 
                           n16716, ZN => n2939);
   U16596 : OAI22_X1 port map( A1 => n17915, A2 => n16717, B1 => n16774, B2 => 
                           n16716, ZN => n2938);
   U16597 : OAI22_X1 port map( A1 => n17916, A2 => n16715, B1 => n16775, B2 => 
                           n16716, ZN => n2937);
   U16598 : OAI22_X1 port map( A1 => n17917, A2 => n16717, B1 => n16776, B2 => 
                           n16716, ZN => n2936);
   U16599 : OAI22_X1 port map( A1 => n17317, A2 => n16715, B1 => n16777, B2 => 
                           n16716, ZN => n2935);
   U16600 : OAI22_X1 port map( A1 => n17318, A2 => n16717, B1 => n16778, B2 => 
                           n16716, ZN => n2934);
   U16601 : OAI22_X1 port map( A1 => n17658, A2 => n16715, B1 => n16779, B2 => 
                           n16716, ZN => n2933);
   U16602 : OAI22_X1 port map( A1 => n17319, A2 => n16717, B1 => n16781, B2 => 
                           n16718, ZN => n2932);
   U16603 : OAI22_X1 port map( A1 => n17018, A2 => n16717, B1 => n16782, B2 => 
                           n16718, ZN => n2931);
   U16604 : OAI22_X1 port map( A1 => n17019, A2 => n16715, B1 => n16783, B2 => 
                           n16718, ZN => n2930);
   U16605 : OAI22_X1 port map( A1 => n17126, A2 => n16717, B1 => n16784, B2 => 
                           n16718, ZN => n2929);
   U16606 : OAI22_X1 port map( A1 => n17127, A2 => n16715, B1 => n16785, B2 => 
                           n16718, ZN => n2928);
   U16607 : OAI22_X1 port map( A1 => n17020, A2 => n16717, B1 => n16786, B2 => 
                           n16718, ZN => n2927);
   U16608 : OAI22_X1 port map( A1 => n16922, A2 => n16715, B1 => n16787, B2 => 
                           n16718, ZN => n2926);
   U16609 : OAI22_X1 port map( A1 => n17021, A2 => n16715, B1 => n16788, B2 => 
                           n16718, ZN => n2925);
   U16610 : OAI22_X1 port map( A1 => n17022, A2 => n16715, B1 => n16789, B2 => 
                           n16718, ZN => n2924);
   U16611 : OAI22_X1 port map( A1 => n16923, A2 => n16715, B1 => n16790, B2 => 
                           n16718, ZN => n2923);
   U16612 : OAI22_X1 port map( A1 => n17023, A2 => n16715, B1 => n16791, B2 => 
                           n16718, ZN => n2922);
   U16613 : OAI22_X1 port map( A1 => n17128, A2 => n16715, B1 => n16792, B2 => 
                           n16718, ZN => n2921);
   U16614 : OAI22_X1 port map( A1 => n17024, A2 => n16715, B1 => n16793, B2 => 
                           n16718, ZN => n2920);
   U16615 : OAI22_X1 port map( A1 => n17320, A2 => n16717, B1 => n16794, B2 => 
                           n16718, ZN => n2919);
   U16616 : OAI22_X1 port map( A1 => n17918, A2 => n16717, B1 => n16795, B2 => 
                           n16718, ZN => n2918);
   U16617 : OAI22_X1 port map( A1 => n17659, A2 => n16715, B1 => n16796, B2 => 
                           n16718, ZN => n2917);
   U16618 : OAI22_X1 port map( A1 => n17660, A2 => n16715, B1 => n16797, B2 => 
                           n16718, ZN => n2916);
   U16619 : OAI22_X1 port map( A1 => n17321, A2 => n16717, B1 => n16798, B2 => 
                           n16718, ZN => n2915);
   U16620 : OAI22_X1 port map( A1 => n17919, A2 => n16715, B1 => n16799, B2 => 
                           n16718, ZN => n2914);
   U16621 : OAI22_X1 port map( A1 => n17322, A2 => n16717, B1 => n16800, B2 => 
                           n16718, ZN => n2913);
   U16622 : OAI22_X1 port map( A1 => n17920, A2 => n16715, B1 => n16801, B2 => 
                           n16718, ZN => n2912);
   U16623 : OAI22_X1 port map( A1 => n17921, A2 => n16717, B1 => n16802, B2 => 
                           n16718, ZN => n2911);
   U16624 : OAI22_X1 port map( A1 => n17661, A2 => n16717, B1 => n16803, B2 => 
                           n16718, ZN => n2910);
   U16625 : OAI22_X1 port map( A1 => n17662, A2 => n16715, B1 => n16804, B2 => 
                           n16718, ZN => n2909);
   U16626 : OAI22_X1 port map( A1 => n17323, A2 => n16715, B1 => n16805, B2 => 
                           n16716, ZN => n2908);
   U16627 : OAI22_X1 port map( A1 => n17663, A2 => n16717, B1 => n16806, B2 => 
                           n16718, ZN => n2907);
   U16628 : OAI22_X1 port map( A1 => n17922, A2 => n16715, B1 => n16808, B2 => 
                           n16718, ZN => n2906);
   U16629 : OAI22_X1 port map( A1 => n17664, A2 => n16717, B1 => n16810, B2 => 
                           n16716, ZN => n2905);
   U16630 : OAI22_X1 port map( A1 => n17665, A2 => n16715, B1 => n16812, B2 => 
                           n16718, ZN => n2904);
   U16631 : NAND2_X1 port map( A1 => n16719, A2 => n16813, ZN => n16722);
   U16632 : NAND2_X1 port map( A1 => n13731, A2 => n16721, ZN => n16723);
   U16633 : OAI22_X1 port map( A1 => n18241, A2 => n16723, B1 => n16815, B2 => 
                           n16722, ZN => n2903);
   U16634 : CLKBUF_X2 port map( A => n16723, Z => n16720);
   U16635 : CLKBUF_X2 port map( A => n16722, Z => n16721);
   U16636 : OAI22_X1 port map( A1 => n17025, A2 => n16720, B1 => n16816, B2 => 
                           n16721, ZN => n2902);
   U16637 : OAI22_X1 port map( A1 => n16924, A2 => n16723, B1 => n16817, B2 => 
                           n16722, ZN => n2901);
   U16638 : OAI22_X1 port map( A1 => n17129, A2 => n16720, B1 => n16818, B2 => 
                           n16722, ZN => n2900);
   U16639 : OAI22_X1 port map( A1 => n17026, A2 => n16720, B1 => n16819, B2 => 
                           n16722, ZN => n2899);
   U16640 : OAI22_X1 port map( A1 => n17130, A2 => n16720, B1 => n16820, B2 => 
                           n16722, ZN => n2898);
   U16641 : OAI22_X1 port map( A1 => n17027, A2 => n16720, B1 => n16821, B2 => 
                           n16721, ZN => n2897);
   U16642 : OAI22_X1 port map( A1 => n16925, A2 => n16720, B1 => n16822, B2 => 
                           n16722, ZN => n2896);
   U16643 : OAI22_X1 port map( A1 => n17131, A2 => n16720, B1 => n16823, B2 => 
                           n16721, ZN => n2895);
   U16644 : OAI22_X1 port map( A1 => n17132, A2 => n16720, B1 => n16824, B2 => 
                           n16722, ZN => n2894);
   U16645 : OAI22_X1 port map( A1 => n17028, A2 => n16720, B1 => n16825, B2 => 
                           n16721, ZN => n2893);
   U16646 : OAI22_X1 port map( A1 => n17029, A2 => n16720, B1 => n16826, B2 => 
                           n16721, ZN => n2892);
   U16647 : OAI22_X1 port map( A1 => n17666, A2 => n16723, B1 => n16827, B2 => 
                           n16722, ZN => n2891);
   U16648 : OAI22_X1 port map( A1 => n17923, A2 => n16720, B1 => n16828, B2 => 
                           n16721, ZN => n2890);
   U16649 : OAI22_X1 port map( A1 => n17924, A2 => n16720, B1 => n16829, B2 => 
                           n16722, ZN => n2889);
   U16650 : OAI22_X1 port map( A1 => n17925, A2 => n16723, B1 => n16830, B2 => 
                           n16721, ZN => n2888);
   U16651 : OAI22_X1 port map( A1 => n17667, A2 => n16723, B1 => n16831, B2 => 
                           n16722, ZN => n2887);
   U16652 : OAI22_X1 port map( A1 => n17926, A2 => n16720, B1 => n16832, B2 => 
                           n16721, ZN => n2886);
   U16653 : OAI22_X1 port map( A1 => n17927, A2 => n16720, B1 => n16833, B2 => 
                           n16722, ZN => n2885);
   U16654 : OAI22_X1 port map( A1 => n17928, A2 => n16723, B1 => n16834, B2 => 
                           n16721, ZN => n2884);
   U16655 : OAI22_X1 port map( A1 => n17668, A2 => n16723, B1 => n16835, B2 => 
                           n16721, ZN => n2883);
   U16656 : OAI22_X1 port map( A1 => n17669, A2 => n16720, B1 => n16836, B2 => 
                           n16721, ZN => n2882);
   U16657 : OAI22_X1 port map( A1 => n17670, A2 => n16720, B1 => n16837, B2 => 
                           n16721, ZN => n2881);
   U16658 : OAI22_X1 port map( A1 => n17671, A2 => n16720, B1 => n16838, B2 => 
                           n16722, ZN => n2880);
   U16659 : OAI22_X1 port map( A1 => n17324, A2 => n16720, B1 => n16839, B2 => 
                           n16721, ZN => n2879);
   U16660 : OAI22_X1 port map( A1 => n17929, A2 => n16723, B1 => n16840, B2 => 
                           n16722, ZN => n2878);
   U16661 : OAI22_X1 port map( A1 => n17672, A2 => n16720, B1 => n16841, B2 => 
                           n16722, ZN => n2877);
   U16662 : OAI22_X1 port map( A1 => n17930, A2 => n16723, B1 => n16842, B2 => 
                           n16722, ZN => n2876);
   U16663 : OAI22_X1 port map( A1 => n17931, A2 => n16720, B1 => n16843, B2 => 
                           n16722, ZN => n2875);
   U16664 : OAI22_X1 port map( A1 => n17673, A2 => n16723, B1 => n16844, B2 => 
                           n16722, ZN => n2874);
   U16665 : OAI22_X1 port map( A1 => n17674, A2 => n16720, B1 => n16845, B2 => 
                           n16722, ZN => n2873);
   U16666 : OAI22_X1 port map( A1 => n17675, A2 => n16723, B1 => n16846, B2 => 
                           n16722, ZN => n2872);
   U16667 : OAI22_X1 port map( A1 => n17676, A2 => n16720, B1 => n16847, B2 => 
                           n16722, ZN => n2871);
   U16668 : OAI22_X1 port map( A1 => n17932, A2 => n16723, B1 => n16848, B2 => 
                           n16722, ZN => n2870);
   U16669 : OAI22_X1 port map( A1 => n17933, A2 => n16720, B1 => n16849, B2 => 
                           n16722, ZN => n2869);
   U16670 : OAI22_X1 port map( A1 => n17934, A2 => n16723, B1 => n16850, B2 => 
                           n16721, ZN => n2868);
   U16671 : OAI22_X1 port map( A1 => n17133, A2 => n16723, B1 => n16851, B2 => 
                           n16721, ZN => n2867);
   U16672 : OAI22_X1 port map( A1 => n17134, A2 => n16720, B1 => n16852, B2 => 
                           n16721, ZN => n2866);
   U16673 : OAI22_X1 port map( A1 => n17030, A2 => n16723, B1 => n16853, B2 => 
                           n16721, ZN => n2865);
   U16674 : OAI22_X1 port map( A1 => n17031, A2 => n16720, B1 => n16854, B2 => 
                           n16721, ZN => n2864);
   U16675 : OAI22_X1 port map( A1 => n17032, A2 => n16723, B1 => n16855, B2 => 
                           n16721, ZN => n2863);
   U16676 : OAI22_X1 port map( A1 => n17033, A2 => n16720, B1 => n16856, B2 => 
                           n16721, ZN => n2862);
   U16677 : OAI22_X1 port map( A1 => n17135, A2 => n16720, B1 => n16857, B2 => 
                           n16721, ZN => n2861);
   U16678 : OAI22_X1 port map( A1 => n17136, A2 => n16720, B1 => n16858, B2 => 
                           n16721, ZN => n2860);
   U16679 : OAI22_X1 port map( A1 => n16926, A2 => n16720, B1 => n16859, B2 => 
                           n16721, ZN => n2859);
   U16680 : OAI22_X1 port map( A1 => n17034, A2 => n16720, B1 => n16860, B2 => 
                           n16721, ZN => n2858);
   U16681 : OAI22_X1 port map( A1 => n17137, A2 => n16720, B1 => n16861, B2 => 
                           n16721, ZN => n2857);
   U16682 : OAI22_X1 port map( A1 => n16927, A2 => n16720, B1 => n16862, B2 => 
                           n16721, ZN => n2856);
   U16683 : OAI22_X1 port map( A1 => n17677, A2 => n16723, B1 => n16863, B2 => 
                           n16721, ZN => n2855);
   U16684 : OAI22_X1 port map( A1 => n17678, A2 => n16723, B1 => n16864, B2 => 
                           n16721, ZN => n2854);
   U16685 : OAI22_X1 port map( A1 => n17679, A2 => n16720, B1 => n16865, B2 => 
                           n16721, ZN => n2853);
   U16686 : OAI22_X1 port map( A1 => n17680, A2 => n16720, B1 => n16866, B2 => 
                           n16721, ZN => n2852);
   U16687 : OAI22_X1 port map( A1 => n17325, A2 => n16723, B1 => n16867, B2 => 
                           n16721, ZN => n2851);
   U16688 : OAI22_X1 port map( A1 => n17681, A2 => n16720, B1 => n16868, B2 => 
                           n16721, ZN => n2850);
   U16689 : OAI22_X1 port map( A1 => n17682, A2 => n16723, B1 => n16869, B2 => 
                           n16721, ZN => n2849);
   U16690 : OAI22_X1 port map( A1 => n17683, A2 => n16720, B1 => n16870, B2 => 
                           n16721, ZN => n2848);
   U16691 : OAI22_X1 port map( A1 => n17684, A2 => n16723, B1 => n16871, B2 => 
                           n16721, ZN => n2847);
   U16692 : OAI22_X1 port map( A1 => n17935, A2 => n16723, B1 => n16872, B2 => 
                           n16721, ZN => n2846);
   U16693 : OAI22_X1 port map( A1 => n17936, A2 => n16720, B1 => n16873, B2 => 
                           n16721, ZN => n2845);
   U16694 : OAI22_X1 port map( A1 => n17937, A2 => n16720, B1 => n16874, B2 => 
                           n16722, ZN => n2844);
   U16695 : OAI22_X1 port map( A1 => n17938, A2 => n16723, B1 => n16875, B2 => 
                           n16721, ZN => n2843);
   U16696 : OAI22_X1 port map( A1 => n17939, A2 => n16720, B1 => n16876, B2 => 
                           n16721, ZN => n2842);
   U16697 : OAI22_X1 port map( A1 => n17940, A2 => n16723, B1 => n16878, B2 => 
                           n16722, ZN => n2841);
   U16698 : OAI22_X1 port map( A1 => n17685, A2 => n16720, B1 => n16881, B2 => 
                           n16721, ZN => n2840);
   U16699 : NAND2_X1 port map( A1 => n16724, A2 => n16813, ZN => n16726);
   U16700 : CLKBUF_X2 port map( A => n16726, Z => n16728);
   U16701 : NAND2_X1 port map( A1 => n13731, A2 => n16728, ZN => n16727);
   U16702 : OAI22_X1 port map( A1 => n18699, A2 => n16727, B1 => n16745, B2 => 
                           n16726, ZN => n2839);
   U16703 : CLKBUF_X2 port map( A => n16727, Z => n16725);
   U16704 : OAI22_X1 port map( A1 => n17138, A2 => n16725, B1 => n16746, B2 => 
                           n16728, ZN => n2838);
   U16705 : OAI22_X1 port map( A1 => n17035, A2 => n16727, B1 => n16747, B2 => 
                           n16726, ZN => n2837);
   U16706 : OAI22_X1 port map( A1 => n17036, A2 => n16725, B1 => n16748, B2 => 
                           n16726, ZN => n2836);
   U16707 : OAI22_X1 port map( A1 => n17139, A2 => n16725, B1 => n16749, B2 => 
                           n16728, ZN => n2835);
   U16708 : OAI22_X1 port map( A1 => n17037, A2 => n16725, B1 => n16750, B2 => 
                           n16726, ZN => n2834);
   U16709 : OAI22_X1 port map( A1 => n17038, A2 => n16725, B1 => n16751, B2 => 
                           n16728, ZN => n2833);
   U16710 : OAI22_X1 port map( A1 => n17140, A2 => n16725, B1 => n16752, B2 => 
                           n16728, ZN => n2832);
   U16711 : OAI22_X1 port map( A1 => n17141, A2 => n16725, B1 => n16753, B2 => 
                           n16728, ZN => n2831);
   U16712 : OAI22_X1 port map( A1 => n17039, A2 => n16725, B1 => n16754, B2 => 
                           n16728, ZN => n2830);
   U16713 : OAI22_X1 port map( A1 => n17142, A2 => n16725, B1 => n16755, B2 => 
                           n16728, ZN => n2829);
   U16714 : OAI22_X1 port map( A1 => n17143, A2 => n16725, B1 => n16756, B2 => 
                           n16726, ZN => n2828);
   U16715 : OAI22_X1 port map( A1 => n17941, A2 => n16727, B1 => n16757, B2 => 
                           n16726, ZN => n2827);
   U16716 : OAI22_X1 port map( A1 => n17942, A2 => n16725, B1 => n16758, B2 => 
                           n16728, ZN => n2826);
   U16717 : OAI22_X1 port map( A1 => n17943, A2 => n16725, B1 => n16759, B2 => 
                           n16726, ZN => n2825);
   U16718 : OAI22_X1 port map( A1 => n17686, A2 => n16727, B1 => n16760, B2 => 
                           n16726, ZN => n2824);
   U16719 : OAI22_X1 port map( A1 => n17944, A2 => n16727, B1 => n16761, B2 => 
                           n16726, ZN => n2823);
   U16720 : OAI22_X1 port map( A1 => n17687, A2 => n16725, B1 => n16762, B2 => 
                           n16728, ZN => n2822);
   U16721 : OAI22_X1 port map( A1 => n17688, A2 => n16725, B1 => n16763, B2 => 
                           n16726, ZN => n2821);
   U16722 : OAI22_X1 port map( A1 => n17945, A2 => n16727, B1 => n16764, B2 => 
                           n16726, ZN => n2820);
   U16723 : OAI22_X1 port map( A1 => n17689, A2 => n16727, B1 => n16765, B2 => 
                           n16728, ZN => n2819);
   U16724 : OAI22_X1 port map( A1 => n17946, A2 => n16725, B1 => n16766, B2 => 
                           n16728, ZN => n2818);
   U16725 : OAI22_X1 port map( A1 => n17690, A2 => n16725, B1 => n16767, B2 => 
                           n16728, ZN => n2817);
   U16726 : OAI22_X1 port map( A1 => n17691, A2 => n16725, B1 => n16768, B2 => 
                           n16726, ZN => n2816);
   U16727 : OAI22_X1 port map( A1 => n17692, A2 => n16725, B1 => n16769, B2 => 
                           n16728, ZN => n2815);
   U16728 : OAI22_X1 port map( A1 => n17947, A2 => n16727, B1 => n16770, B2 => 
                           n16726, ZN => n2814);
   U16729 : OAI22_X1 port map( A1 => n17948, A2 => n16725, B1 => n16771, B2 => 
                           n16726, ZN => n2813);
   U16730 : OAI22_X1 port map( A1 => n17949, A2 => n16727, B1 => n16772, B2 => 
                           n16726, ZN => n2812);
   U16731 : OAI22_X1 port map( A1 => n17950, A2 => n16725, B1 => n16773, B2 => 
                           n16726, ZN => n2811);
   U16732 : OAI22_X1 port map( A1 => n17951, A2 => n16727, B1 => n16774, B2 => 
                           n16726, ZN => n2810);
   U16733 : OAI22_X1 port map( A1 => n17693, A2 => n16725, B1 => n16775, B2 => 
                           n16726, ZN => n2809);
   U16734 : OAI22_X1 port map( A1 => n17694, A2 => n16727, B1 => n16776, B2 => 
                           n16726, ZN => n2808);
   U16735 : OAI22_X1 port map( A1 => n17695, A2 => n16725, B1 => n16777, B2 => 
                           n16726, ZN => n2807);
   U16736 : OAI22_X1 port map( A1 => n17696, A2 => n16727, B1 => n16778, B2 => 
                           n16726, ZN => n2806);
   U16737 : OAI22_X1 port map( A1 => n17952, A2 => n16725, B1 => n16779, B2 => 
                           n16726, ZN => n2805);
   U16738 : OAI22_X1 port map( A1 => n17953, A2 => n16727, B1 => n16781, B2 => 
                           n16728, ZN => n2804);
   U16739 : OAI22_X1 port map( A1 => n17040, A2 => n16727, B1 => n16782, B2 => 
                           n16728, ZN => n2803);
   U16740 : OAI22_X1 port map( A1 => n17144, A2 => n16725, B1 => n16783, B2 => 
                           n16728, ZN => n2802);
   U16741 : OAI22_X1 port map( A1 => n17145, A2 => n16727, B1 => n16784, B2 => 
                           n16728, ZN => n2801);
   U16742 : OAI22_X1 port map( A1 => n17041, A2 => n16725, B1 => n16785, B2 => 
                           n16728, ZN => n2800);
   U16743 : OAI22_X1 port map( A1 => n17042, A2 => n16727, B1 => n16786, B2 => 
                           n16728, ZN => n2799);
   U16744 : OAI22_X1 port map( A1 => n17146, A2 => n16725, B1 => n16787, B2 => 
                           n16728, ZN => n2798);
   U16745 : OAI22_X1 port map( A1 => n17147, A2 => n16725, B1 => n16788, B2 => 
                           n16728, ZN => n2797);
   U16746 : OAI22_X1 port map( A1 => n17043, A2 => n16725, B1 => n16789, B2 => 
                           n16728, ZN => n2796);
   U16747 : OAI22_X1 port map( A1 => n17044, A2 => n16725, B1 => n16790, B2 => 
                           n16728, ZN => n2795);
   U16748 : OAI22_X1 port map( A1 => n17045, A2 => n16725, B1 => n16791, B2 => 
                           n16728, ZN => n2794);
   U16749 : OAI22_X1 port map( A1 => n17148, A2 => n16725, B1 => n16792, B2 => 
                           n16728, ZN => n2793);
   U16750 : OAI22_X1 port map( A1 => n17149, A2 => n16725, B1 => n16793, B2 => 
                           n16728, ZN => n2792);
   U16751 : OAI22_X1 port map( A1 => n17954, A2 => n16727, B1 => n16794, B2 => 
                           n16728, ZN => n2791);
   U16752 : OAI22_X1 port map( A1 => n17955, A2 => n16727, B1 => n16795, B2 => 
                           n16728, ZN => n2790);
   U16753 : OAI22_X1 port map( A1 => n17956, A2 => n16725, B1 => n16796, B2 => 
                           n16728, ZN => n2789);
   U16754 : OAI22_X1 port map( A1 => n17697, A2 => n16725, B1 => n16797, B2 => 
                           n16728, ZN => n2788);
   U16755 : OAI22_X1 port map( A1 => n17957, A2 => n16727, B1 => n16798, B2 => 
                           n16728, ZN => n2787);
   U16756 : OAI22_X1 port map( A1 => n17698, A2 => n16725, B1 => n16799, B2 => 
                           n16728, ZN => n2786);
   U16757 : OAI22_X1 port map( A1 => n17958, A2 => n16727, B1 => n16800, B2 => 
                           n16728, ZN => n2785);
   U16758 : OAI22_X1 port map( A1 => n17959, A2 => n16725, B1 => n16801, B2 => 
                           n16728, ZN => n2784);
   U16759 : OAI22_X1 port map( A1 => n17699, A2 => n16727, B1 => n16802, B2 => 
                           n16728, ZN => n2783);
   U16760 : OAI22_X1 port map( A1 => n17700, A2 => n16727, B1 => n16803, B2 => 
                           n16728, ZN => n2782);
   U16761 : OAI22_X1 port map( A1 => n17701, A2 => n16725, B1 => n16804, B2 => 
                           n16728, ZN => n2781);
   U16762 : OAI22_X1 port map( A1 => n17960, A2 => n16725, B1 => n16805, B2 => 
                           n16726, ZN => n2780);
   U16763 : OAI22_X1 port map( A1 => n17961, A2 => n16727, B1 => n16806, B2 => 
                           n16728, ZN => n2779);
   U16764 : OAI22_X1 port map( A1 => n17962, A2 => n16725, B1 => n16808, B2 => 
                           n16728, ZN => n2778);
   U16765 : OAI22_X1 port map( A1 => n17702, A2 => n16727, B1 => n16810, B2 => 
                           n16726, ZN => n2777);
   U16766 : OAI22_X1 port map( A1 => n17703, A2 => n16725, B1 => n16812, B2 => 
                           n16728, ZN => n2776);
   U16767 : NAND2_X1 port map( A1 => n16729, A2 => n16813, ZN => n16731);
   U16768 : CLKBUF_X2 port map( A => n16731, Z => n16733);
   U16769 : NAND2_X1 port map( A1 => n13731, A2 => n16733, ZN => n16732);
   U16770 : OAI22_X1 port map( A1 => n18014, A2 => n16732, B1 => n16815, B2 => 
                           n16731, ZN => n2775);
   U16771 : CLKBUF_X2 port map( A => n16732, Z => n16730);
   U16772 : OAI22_X1 port map( A1 => n17150, A2 => n16730, B1 => n16816, B2 => 
                           n16733, ZN => n2774);
   U16773 : OAI22_X1 port map( A1 => n16928, A2 => n16732, B1 => n16817, B2 => 
                           n16731, ZN => n2773);
   U16774 : OAI22_X1 port map( A1 => n17046, A2 => n16730, B1 => n16818, B2 => 
                           n16731, ZN => n2772);
   U16775 : OAI22_X1 port map( A1 => n17151, A2 => n16730, B1 => n16819, B2 => 
                           n16733, ZN => n2771);
   U16776 : OAI22_X1 port map( A1 => n17047, A2 => n16730, B1 => n16820, B2 => 
                           n16731, ZN => n2770);
   U16777 : OAI22_X1 port map( A1 => n16929, A2 => n16730, B1 => n16821, B2 => 
                           n16733, ZN => n2769);
   U16778 : OAI22_X1 port map( A1 => n17152, A2 => n16730, B1 => n16822, B2 => 
                           n16733, ZN => n2768);
   U16779 : OAI22_X1 port map( A1 => n16930, A2 => n16730, B1 => n16823, B2 => 
                           n16733, ZN => n2767);
   U16780 : OAI22_X1 port map( A1 => n17048, A2 => n16730, B1 => n16824, B2 => 
                           n16733, ZN => n2766);
   U16781 : OAI22_X1 port map( A1 => n17049, A2 => n16730, B1 => n16825, B2 => 
                           n16733, ZN => n2765);
   U16782 : OAI22_X1 port map( A1 => n17050, A2 => n16730, B1 => n16826, B2 => 
                           n16731, ZN => n2764);
   U16783 : OAI22_X1 port map( A1 => n17326, A2 => n16732, B1 => n16827, B2 => 
                           n16731, ZN => n2763);
   U16784 : OAI22_X1 port map( A1 => n17963, A2 => n16730, B1 => n16828, B2 => 
                           n16733, ZN => n2762);
   U16785 : OAI22_X1 port map( A1 => n17704, A2 => n16730, B1 => n16829, B2 => 
                           n16731, ZN => n2761);
   U16786 : OAI22_X1 port map( A1 => n17705, A2 => n16732, B1 => n16830, B2 => 
                           n16731, ZN => n2760);
   U16787 : OAI22_X1 port map( A1 => n17964, A2 => n16732, B1 => n16831, B2 => 
                           n16731, ZN => n2759);
   U16788 : OAI22_X1 port map( A1 => n17706, A2 => n16730, B1 => n16832, B2 => 
                           n16733, ZN => n2758);
   U16789 : OAI22_X1 port map( A1 => n17327, A2 => n16730, B1 => n16833, B2 => 
                           n16731, ZN => n2757);
   U16790 : OAI22_X1 port map( A1 => n17965, A2 => n16732, B1 => n16834, B2 => 
                           n16731, ZN => n2756);
   U16791 : OAI22_X1 port map( A1 => n17328, A2 => n16732, B1 => n16835, B2 => 
                           n16733, ZN => n2755);
   U16792 : OAI22_X1 port map( A1 => n17707, A2 => n16730, B1 => n16836, B2 => 
                           n16733, ZN => n2754);
   U16793 : OAI22_X1 port map( A1 => n17966, A2 => n16730, B1 => n16837, B2 => 
                           n16733, ZN => n2753);
   U16794 : OAI22_X1 port map( A1 => n17967, A2 => n16730, B1 => n16838, B2 => 
                           n16731, ZN => n2752);
   U16795 : OAI22_X1 port map( A1 => n17968, A2 => n16730, B1 => n16839, B2 => 
                           n16733, ZN => n2751);
   U16796 : OAI22_X1 port map( A1 => n17708, A2 => n16732, B1 => n16840, B2 => 
                           n16731, ZN => n2750);
   U16797 : OAI22_X1 port map( A1 => n17969, A2 => n16730, B1 => n16841, B2 => 
                           n16731, ZN => n2749);
   U16798 : OAI22_X1 port map( A1 => n17709, A2 => n16732, B1 => n16842, B2 => 
                           n16731, ZN => n2748);
   U16799 : OAI22_X1 port map( A1 => n17970, A2 => n16730, B1 => n16843, B2 => 
                           n16731, ZN => n2747);
   U16800 : OAI22_X1 port map( A1 => n17710, A2 => n16732, B1 => n16844, B2 => 
                           n16731, ZN => n2746);
   U16801 : OAI22_X1 port map( A1 => n17711, A2 => n16730, B1 => n16845, B2 => 
                           n16731, ZN => n2745);
   U16802 : OAI22_X1 port map( A1 => n17971, A2 => n16732, B1 => n16846, B2 => 
                           n16731, ZN => n2744);
   U16803 : OAI22_X1 port map( A1 => n17972, A2 => n16730, B1 => n16847, B2 => 
                           n16731, ZN => n2743);
   U16804 : OAI22_X1 port map( A1 => n17712, A2 => n16732, B1 => n16848, B2 => 
                           n16731, ZN => n2742);
   U16805 : OAI22_X1 port map( A1 => n17713, A2 => n16730, B1 => n16849, B2 => 
                           n16731, ZN => n2741);
   U16806 : OAI22_X1 port map( A1 => n17714, A2 => n16732, B1 => n16850, B2 => 
                           n16733, ZN => n2740);
   U16807 : OAI22_X1 port map( A1 => n17153, A2 => n16732, B1 => n16851, B2 => 
                           n16733, ZN => n2739);
   U16808 : OAI22_X1 port map( A1 => n17154, A2 => n16730, B1 => n16852, B2 => 
                           n16733, ZN => n2738);
   U16809 : OAI22_X1 port map( A1 => n17155, A2 => n16732, B1 => n16853, B2 => 
                           n16733, ZN => n2737);
   U16810 : OAI22_X1 port map( A1 => n17156, A2 => n16730, B1 => n16854, B2 => 
                           n16733, ZN => n2736);
   U16811 : OAI22_X1 port map( A1 => n17051, A2 => n16732, B1 => n16855, B2 => 
                           n16733, ZN => n2735);
   U16812 : OAI22_X1 port map( A1 => n17052, A2 => n16730, B1 => n16856, B2 => 
                           n16733, ZN => n2734);
   U16813 : OAI22_X1 port map( A1 => n16931, A2 => n16730, B1 => n16857, B2 => 
                           n16733, ZN => n2733);
   U16814 : OAI22_X1 port map( A1 => n17053, A2 => n16730, B1 => n16858, B2 => 
                           n16733, ZN => n2732);
   U16815 : OAI22_X1 port map( A1 => n17157, A2 => n16730, B1 => n16859, B2 => 
                           n16733, ZN => n2731);
   U16816 : OAI22_X1 port map( A1 => n17158, A2 => n16730, B1 => n16860, B2 => 
                           n16733, ZN => n2730);
   U16817 : OAI22_X1 port map( A1 => n17054, A2 => n16730, B1 => n16861, B2 => 
                           n16733, ZN => n2729);
   U16818 : OAI22_X1 port map( A1 => n16932, A2 => n16730, B1 => n16862, B2 => 
                           n16733, ZN => n2728);
   U16819 : OAI22_X1 port map( A1 => n17973, A2 => n16732, B1 => n16863, B2 => 
                           n16733, ZN => n2727);
   U16820 : OAI22_X1 port map( A1 => n17329, A2 => n16732, B1 => n16864, B2 => 
                           n16733, ZN => n2726);
   U16821 : OAI22_X1 port map( A1 => n17715, A2 => n16730, B1 => n16865, B2 => 
                           n16733, ZN => n2725);
   U16822 : OAI22_X1 port map( A1 => n17974, A2 => n16730, B1 => n16866, B2 => 
                           n16733, ZN => n2724);
   U16823 : OAI22_X1 port map( A1 => n17716, A2 => n16732, B1 => n16867, B2 => 
                           n16733, ZN => n2723);
   U16824 : OAI22_X1 port map( A1 => n17975, A2 => n16730, B1 => n16868, B2 => 
                           n16733, ZN => n2722);
   U16825 : OAI22_X1 port map( A1 => n17717, A2 => n16732, B1 => n16869, B2 => 
                           n16733, ZN => n2721);
   U16826 : OAI22_X1 port map( A1 => n17718, A2 => n16730, B1 => n16870, B2 => 
                           n16733, ZN => n2720);
   U16827 : OAI22_X1 port map( A1 => n17976, A2 => n16732, B1 => n16871, B2 => 
                           n16733, ZN => n2719);
   U16828 : OAI22_X1 port map( A1 => n17977, A2 => n16732, B1 => n16872, B2 => 
                           n16733, ZN => n2718);
   U16829 : OAI22_X1 port map( A1 => n17719, A2 => n16730, B1 => n16873, B2 => 
                           n16733, ZN => n2717);
   U16830 : OAI22_X1 port map( A1 => n17720, A2 => n16730, B1 => n16874, B2 => 
                           n16731, ZN => n2716);
   U16831 : OAI22_X1 port map( A1 => n17721, A2 => n16732, B1 => n16875, B2 => 
                           n16733, ZN => n2715);
   U16832 : OAI22_X1 port map( A1 => n17330, A2 => n16730, B1 => n16876, B2 => 
                           n16733, ZN => n2714);
   U16833 : OAI22_X1 port map( A1 => n17978, A2 => n16732, B1 => n16878, B2 => 
                           n16731, ZN => n2713);
   U16834 : OAI22_X1 port map( A1 => n17722, A2 => n16730, B1 => n16881, B2 => 
                           n16733, ZN => n2712);
   U16835 : NAND2_X1 port map( A1 => n16734, A2 => n16813, ZN => n16735);
   U16836 : CLKBUF_X2 port map( A => n16735, Z => n16737);
   U16837 : NAND2_X1 port map( A1 => n13731, A2 => n16737, ZN => n16736);
   U16838 : OAI22_X1 port map( A1 => n18700, A2 => n16736, B1 => n16745, B2 => 
                           n16735, ZN => n2711);
   U16839 : OAI22_X1 port map( A1 => n16933, A2 => n16738, B1 => n16746, B2 => 
                           n16737, ZN => n2710);
   U16840 : OAI22_X1 port map( A1 => n17055, A2 => n16736, B1 => n16747, B2 => 
                           n16735, ZN => n2709);
   U16841 : OAI22_X1 port map( A1 => n16934, A2 => n16738, B1 => n16748, B2 => 
                           n16735, ZN => n2708);
   U16842 : OAI22_X1 port map( A1 => n17056, A2 => n16738, B1 => n16749, B2 => 
                           n16737, ZN => n2707);
   U16843 : OAI22_X1 port map( A1 => n17057, A2 => n16736, B1 => n16750, B2 => 
                           n16735, ZN => n2706);
   U16844 : OAI22_X1 port map( A1 => n17058, A2 => n16738, B1 => n16751, B2 => 
                           n16737, ZN => n2705);
   U16845 : OAI22_X1 port map( A1 => n17059, A2 => n16736, B1 => n16752, B2 => 
                           n16737, ZN => n2704);
   U16846 : OAI22_X1 port map( A1 => n17060, A2 => n16738, B1 => n16753, B2 => 
                           n16737, ZN => n2703);
   U16847 : OAI22_X1 port map( A1 => n17061, A2 => n16736, B1 => n16754, B2 => 
                           n16737, ZN => n2702);
   U16848 : OAI22_X1 port map( A1 => n17062, A2 => n16738, B1 => n16755, B2 => 
                           n16737, ZN => n2701);
   U16849 : OAI22_X1 port map( A1 => n16935, A2 => n16738, B1 => n16756, B2 => 
                           n16735, ZN => n2700);
   U16850 : OAI22_X1 port map( A1 => n17723, A2 => n16736, B1 => n16757, B2 => 
                           n16735, ZN => n2699);
   U16851 : OAI22_X1 port map( A1 => n17724, A2 => n16738, B1 => n16758, B2 => 
                           n16737, ZN => n2698);
   U16852 : OAI22_X1 port map( A1 => n17725, A2 => n16738, B1 => n16759, B2 => 
                           n16735, ZN => n2697);
   U16853 : OAI22_X1 port map( A1 => n17979, A2 => n16736, B1 => n16760, B2 => 
                           n16735, ZN => n2696);
   U16854 : OAI22_X1 port map( A1 => n17331, A2 => n16736, B1 => n16761, B2 => 
                           n16735, ZN => n2695);
   U16855 : OAI22_X1 port map( A1 => n17726, A2 => n16738, B1 => n16762, B2 => 
                           n16737, ZN => n2694);
   U16856 : OAI22_X1 port map( A1 => n17727, A2 => n16738, B1 => n16763, B2 => 
                           n16735, ZN => n2693);
   U16857 : OAI22_X1 port map( A1 => n17728, A2 => n16736, B1 => n16764, B2 => 
                           n16735, ZN => n2692);
   U16858 : OAI22_X1 port map( A1 => n17729, A2 => n16736, B1 => n16765, B2 => 
                           n16737, ZN => n2691);
   U16859 : OAI22_X1 port map( A1 => n17332, A2 => n16738, B1 => n16766, B2 => 
                           n16737, ZN => n2690);
   U16860 : OAI22_X1 port map( A1 => n17333, A2 => n16738, B1 => n16767, B2 => 
                           n16737, ZN => n2689);
   U16861 : OAI22_X1 port map( A1 => n17334, A2 => n16738, B1 => n16768, B2 => 
                           n16735, ZN => n2688);
   U16862 : OAI22_X1 port map( A1 => n17335, A2 => n16738, B1 => n16769, B2 => 
                           n16737, ZN => n2687);
   U16863 : OAI22_X1 port map( A1 => n17730, A2 => n16736, B1 => n16770, B2 => 
                           n16735, ZN => n2686);
   U16864 : OAI22_X1 port map( A1 => n17731, A2 => n16738, B1 => n16771, B2 => 
                           n16735, ZN => n2685);
   U16865 : OAI22_X1 port map( A1 => n17732, A2 => n16736, B1 => n16772, B2 => 
                           n16735, ZN => n2684);
   U16866 : OAI22_X1 port map( A1 => n17336, A2 => n16738, B1 => n16773, B2 => 
                           n16735, ZN => n2683);
   U16867 : OAI22_X1 port map( A1 => n17733, A2 => n16736, B1 => n16774, B2 => 
                           n16735, ZN => n2682);
   U16868 : OAI22_X1 port map( A1 => n17734, A2 => n16738, B1 => n16775, B2 => 
                           n16735, ZN => n2681);
   U16869 : OAI22_X1 port map( A1 => n17735, A2 => n16736, B1 => n16776, B2 => 
                           n16735, ZN => n2680);
   U16870 : OAI22_X1 port map( A1 => n17736, A2 => n16738, B1 => n16777, B2 => 
                           n16735, ZN => n2679);
   U16871 : OAI22_X1 port map( A1 => n17980, A2 => n16736, B1 => n16778, B2 => 
                           n16735, ZN => n2678);
   U16872 : OAI22_X1 port map( A1 => n17337, A2 => n16738, B1 => n16779, B2 => 
                           n16735, ZN => n2677);
   U16873 : OAI22_X1 port map( A1 => n17737, A2 => n16736, B1 => n16781, B2 => 
                           n16737, ZN => n2676);
   U16874 : CLKBUF_X2 port map( A => n16736, Z => n16738);
   U16875 : OAI22_X1 port map( A1 => n17063, A2 => n16738, B1 => n16782, B2 => 
                           n16737, ZN => n2675);
   U16876 : OAI22_X1 port map( A1 => n16936, A2 => n16738, B1 => n16783, B2 => 
                           n16737, ZN => n2674);
   U16877 : OAI22_X1 port map( A1 => n16937, A2 => n16738, B1 => n16784, B2 => 
                           n16737, ZN => n2673);
   U16878 : OAI22_X1 port map( A1 => n17064, A2 => n16738, B1 => n16785, B2 => 
                           n16737, ZN => n2672);
   U16879 : OAI22_X1 port map( A1 => n16938, A2 => n16738, B1 => n16786, B2 => 
                           n16737, ZN => n2671);
   U16880 : OAI22_X1 port map( A1 => n17065, A2 => n16738, B1 => n16787, B2 => 
                           n16737, ZN => n2670);
   U16881 : OAI22_X1 port map( A1 => n16939, A2 => n16738, B1 => n16788, B2 => 
                           n16737, ZN => n2669);
   U16882 : OAI22_X1 port map( A1 => n17066, A2 => n16738, B1 => n16789, B2 => 
                           n16737, ZN => n2668);
   U16883 : OAI22_X1 port map( A1 => n17067, A2 => n16738, B1 => n16790, B2 => 
                           n16737, ZN => n2667);
   U16884 : OAI22_X1 port map( A1 => n16940, A2 => n16738, B1 => n16791, B2 => 
                           n16737, ZN => n2666);
   U16885 : OAI22_X1 port map( A1 => n16941, A2 => n16738, B1 => n16792, B2 => 
                           n16737, ZN => n2665);
   U16886 : OAI22_X1 port map( A1 => n17068, A2 => n16738, B1 => n16793, B2 => 
                           n16737, ZN => n2664);
   U16887 : OAI22_X1 port map( A1 => n17981, A2 => n16736, B1 => n16794, B2 => 
                           n16737, ZN => n2663);
   U16888 : OAI22_X1 port map( A1 => n17338, A2 => n16736, B1 => n16795, B2 => 
                           n16737, ZN => n2662);
   U16889 : OAI22_X1 port map( A1 => n17738, A2 => n16738, B1 => n16796, B2 => 
                           n16737, ZN => n2661);
   U16890 : OAI22_X1 port map( A1 => n17739, A2 => n16738, B1 => n16797, B2 => 
                           n16737, ZN => n2660);
   U16891 : OAI22_X1 port map( A1 => n17339, A2 => n16736, B1 => n16798, B2 => 
                           n16737, ZN => n2659);
   U16892 : OAI22_X1 port map( A1 => n17340, A2 => n16738, B1 => n16799, B2 => 
                           n16737, ZN => n2658);
   U16893 : OAI22_X1 port map( A1 => n17740, A2 => n16736, B1 => n16800, B2 => 
                           n16737, ZN => n2657);
   U16894 : OAI22_X1 port map( A1 => n17741, A2 => n16738, B1 => n16801, B2 => 
                           n16737, ZN => n2656);
   U16895 : OAI22_X1 port map( A1 => n17341, A2 => n16736, B1 => n16802, B2 => 
                           n16737, ZN => n2655);
   U16896 : OAI22_X1 port map( A1 => n17742, A2 => n16736, B1 => n16803, B2 => 
                           n16737, ZN => n2654);
   U16897 : OAI22_X1 port map( A1 => n17743, A2 => n16738, B1 => n16804, B2 => 
                           n16737, ZN => n2653);
   U16898 : OAI22_X1 port map( A1 => n17744, A2 => n16738, B1 => n16805, B2 => 
                           n16735, ZN => n2652);
   U16899 : OAI22_X1 port map( A1 => n17745, A2 => n16736, B1 => n16806, B2 => 
                           n16737, ZN => n2651);
   U16900 : OAI22_X1 port map( A1 => n17746, A2 => n16738, B1 => n16808, B2 => 
                           n16737, ZN => n2650);
   U16901 : OAI22_X1 port map( A1 => n17342, A2 => n16736, B1 => n16810, B2 => 
                           n16735, ZN => n2649);
   U16902 : OAI22_X1 port map( A1 => n17982, A2 => n16738, B1 => n16812, B2 => 
                           n16737, ZN => n2648);
   U16903 : NAND2_X1 port map( A1 => n16739, A2 => n16813, ZN => n16741);
   U16904 : CLKBUF_X2 port map( A => n16741, Z => n16743);
   U16905 : NAND2_X1 port map( A1 => n13731, A2 => n16743, ZN => n16742);
   U16906 : OAI22_X1 port map( A1 => n18015, A2 => n16742, B1 => n16815, B2 => 
                           n16741, ZN => n2647);
   U16907 : CLKBUF_X2 port map( A => n16742, Z => n16740);
   U16908 : OAI22_X1 port map( A1 => n17069, A2 => n16740, B1 => n16816, B2 => 
                           n16743, ZN => n2646);
   U16909 : OAI22_X1 port map( A1 => n17070, A2 => n16742, B1 => n16817, B2 => 
                           n16741, ZN => n2645);
   U16910 : OAI22_X1 port map( A1 => n17071, A2 => n16740, B1 => n16818, B2 => 
                           n16741, ZN => n2644);
   U16911 : OAI22_X1 port map( A1 => n16942, A2 => n16740, B1 => n16819, B2 => 
                           n16743, ZN => n2643);
   U16912 : OAI22_X1 port map( A1 => n17072, A2 => n16740, B1 => n16820, B2 => 
                           n16741, ZN => n2642);
   U16913 : OAI22_X1 port map( A1 => n16943, A2 => n16740, B1 => n16821, B2 => 
                           n16743, ZN => n2641);
   U16914 : OAI22_X1 port map( A1 => n16944, A2 => n16740, B1 => n16822, B2 => 
                           n16743, ZN => n2640);
   U16915 : OAI22_X1 port map( A1 => n16945, A2 => n16740, B1 => n16823, B2 => 
                           n16743, ZN => n2639);
   U16916 : OAI22_X1 port map( A1 => n16946, A2 => n16740, B1 => n16824, B2 => 
                           n16743, ZN => n2638);
   U16917 : OAI22_X1 port map( A1 => n16947, A2 => n16740, B1 => n16825, B2 => 
                           n16743, ZN => n2637);
   U16918 : OAI22_X1 port map( A1 => n16948, A2 => n16740, B1 => n16826, B2 => 
                           n16741, ZN => n2636);
   U16919 : OAI22_X1 port map( A1 => n17747, A2 => n16742, B1 => n16827, B2 => 
                           n16741, ZN => n2635);
   U16920 : OAI22_X1 port map( A1 => n17343, A2 => n16740, B1 => n16828, B2 => 
                           n16743, ZN => n2634);
   U16921 : OAI22_X1 port map( A1 => n17344, A2 => n16740, B1 => n16829, B2 => 
                           n16741, ZN => n2633);
   U16922 : OAI22_X1 port map( A1 => n17345, A2 => n16742, B1 => n16830, B2 => 
                           n16741, ZN => n2632);
   U16923 : OAI22_X1 port map( A1 => n17346, A2 => n16742, B1 => n16831, B2 => 
                           n16741, ZN => n2631);
   U16924 : OAI22_X1 port map( A1 => n17347, A2 => n16740, B1 => n16832, B2 => 
                           n16743, ZN => n2630);
   U16925 : OAI22_X1 port map( A1 => n17748, A2 => n16740, B1 => n16833, B2 => 
                           n16741, ZN => n2629);
   U16926 : OAI22_X1 port map( A1 => n17348, A2 => n16742, B1 => n16834, B2 => 
                           n16741, ZN => n2628);
   U16927 : OAI22_X1 port map( A1 => n17349, A2 => n16742, B1 => n16835, B2 => 
                           n16743, ZN => n2627);
   U16928 : OAI22_X1 port map( A1 => n17350, A2 => n16740, B1 => n16836, B2 => 
                           n16743, ZN => n2626);
   U16929 : OAI22_X1 port map( A1 => n17351, A2 => n16740, B1 => n16837, B2 => 
                           n16743, ZN => n2625);
   U16930 : OAI22_X1 port map( A1 => n17983, A2 => n16740, B1 => n16838, B2 => 
                           n16741, ZN => n2624);
   U16931 : OAI22_X1 port map( A1 => n17749, A2 => n16740, B1 => n16839, B2 => 
                           n16743, ZN => n2623);
   U16932 : OAI22_X1 port map( A1 => n17750, A2 => n16742, B1 => n16840, B2 => 
                           n16741, ZN => n2622);
   U16933 : OAI22_X1 port map( A1 => n17751, A2 => n16740, B1 => n16841, B2 => 
                           n16741, ZN => n2621);
   U16934 : OAI22_X1 port map( A1 => n17984, A2 => n16742, B1 => n16842, B2 => 
                           n16741, ZN => n2620);
   U16935 : OAI22_X1 port map( A1 => n17985, A2 => n16740, B1 => n16843, B2 => 
                           n16741, ZN => n2619);
   U16936 : OAI22_X1 port map( A1 => n17752, A2 => n16742, B1 => n16844, B2 => 
                           n16741, ZN => n2618);
   U16937 : OAI22_X1 port map( A1 => n17753, A2 => n16740, B1 => n16845, B2 => 
                           n16741, ZN => n2617);
   U16938 : OAI22_X1 port map( A1 => n17352, A2 => n16742, B1 => n16846, B2 => 
                           n16741, ZN => n2616);
   U16939 : OAI22_X1 port map( A1 => n17754, A2 => n16740, B1 => n16847, B2 => 
                           n16741, ZN => n2615);
   U16940 : OAI22_X1 port map( A1 => n17353, A2 => n16742, B1 => n16848, B2 => 
                           n16741, ZN => n2614);
   U16941 : OAI22_X1 port map( A1 => n17755, A2 => n16740, B1 => n16849, B2 => 
                           n16741, ZN => n2613);
   U16942 : OAI22_X1 port map( A1 => n17354, A2 => n16742, B1 => n16850, B2 => 
                           n16743, ZN => n2612);
   U16943 : OAI22_X1 port map( A1 => n17073, A2 => n16742, B1 => n16851, B2 => 
                           n16743, ZN => n2611);
   U16944 : OAI22_X1 port map( A1 => n17074, A2 => n16740, B1 => n16852, B2 => 
                           n16743, ZN => n2610);
   U16945 : OAI22_X1 port map( A1 => n16949, A2 => n16742, B1 => n16853, B2 => 
                           n16743, ZN => n2609);
   U16946 : OAI22_X1 port map( A1 => n17075, A2 => n16740, B1 => n16854, B2 => 
                           n16743, ZN => n2608);
   U16947 : OAI22_X1 port map( A1 => n16950, A2 => n16742, B1 => n16855, B2 => 
                           n16743, ZN => n2607);
   U16948 : OAI22_X1 port map( A1 => n17076, A2 => n16740, B1 => n16856, B2 => 
                           n16743, ZN => n2606);
   U16949 : OAI22_X1 port map( A1 => n17077, A2 => n16740, B1 => n16857, B2 => 
                           n16743, ZN => n2605);
   U16950 : OAI22_X1 port map( A1 => n17078, A2 => n16740, B1 => n16858, B2 => 
                           n16743, ZN => n2604);
   U16951 : OAI22_X1 port map( A1 => n16951, A2 => n16740, B1 => n16859, B2 => 
                           n16743, ZN => n2603);
   U16952 : OAI22_X1 port map( A1 => n17079, A2 => n16740, B1 => n16860, B2 => 
                           n16743, ZN => n2602);
   U16953 : OAI22_X1 port map( A1 => n16952, A2 => n16740, B1 => n16861, B2 => 
                           n16743, ZN => n2601);
   U16954 : OAI22_X1 port map( A1 => n16953, A2 => n16740, B1 => n16862, B2 => 
                           n16743, ZN => n2600);
   U16955 : OAI22_X1 port map( A1 => n17986, A2 => n16742, B1 => n16863, B2 => 
                           n16743, ZN => n2599);
   U16956 : OAI22_X1 port map( A1 => n17756, A2 => n16742, B1 => n16864, B2 => 
                           n16743, ZN => n2598);
   U16957 : OAI22_X1 port map( A1 => n17355, A2 => n16740, B1 => n16865, B2 => 
                           n16743, ZN => n2597);
   U16958 : OAI22_X1 port map( A1 => n17356, A2 => n16740, B1 => n16866, B2 => 
                           n16743, ZN => n2596);
   U16959 : OAI22_X1 port map( A1 => n17357, A2 => n16742, B1 => n16867, B2 => 
                           n16743, ZN => n2595);
   U16960 : OAI22_X1 port map( A1 => n17987, A2 => n16740, B1 => n16868, B2 => 
                           n16743, ZN => n2594);
   U16961 : OAI22_X1 port map( A1 => n17757, A2 => n16742, B1 => n16869, B2 => 
                           n16743, ZN => n2593);
   U16962 : OAI22_X1 port map( A1 => n17988, A2 => n16740, B1 => n16870, B2 => 
                           n16743, ZN => n2592);
   U16963 : OAI22_X1 port map( A1 => n17358, A2 => n16742, B1 => n16871, B2 => 
                           n16743, ZN => n2591);
   U16964 : OAI22_X1 port map( A1 => n17359, A2 => n16742, B1 => n16872, B2 => 
                           n16743, ZN => n2590);
   U16965 : OAI22_X1 port map( A1 => n17360, A2 => n16740, B1 => n16873, B2 => 
                           n16743, ZN => n2589);
   U16966 : OAI22_X1 port map( A1 => n17361, A2 => n16740, B1 => n16874, B2 => 
                           n16741, ZN => n2588);
   U16967 : OAI22_X1 port map( A1 => n17362, A2 => n16742, B1 => n16875, B2 => 
                           n16743, ZN => n2587);
   U16968 : OAI22_X1 port map( A1 => n17363, A2 => n16740, B1 => n16876, B2 => 
                           n16743, ZN => n2586);
   U16969 : OAI22_X1 port map( A1 => n17758, A2 => n16742, B1 => n16878, B2 => 
                           n16741, ZN => n2585);
   U16970 : OAI22_X1 port map( A1 => n17759, A2 => n16740, B1 => n16881, B2 => 
                           n16743, ZN => n2584);
   U16971 : NAND2_X1 port map( A1 => n16744, A2 => n16813, ZN => n16809);
   U16972 : NAND2_X1 port map( A1 => n13731, A2 => n16807, ZN => n16811);
   U16973 : OAI22_X1 port map( A1 => n18016, A2 => n16811, B1 => n16745, B2 => 
                           n16809, ZN => n2583);
   U16974 : CLKBUF_X2 port map( A => n16811, Z => n16780);
   U16975 : CLKBUF_X2 port map( A => n16809, Z => n16807);
   U16976 : OAI22_X1 port map( A1 => n17080, A2 => n16780, B1 => n16746, B2 => 
                           n16807, ZN => n2582);
   U16977 : OAI22_X1 port map( A1 => n17081, A2 => n16811, B1 => n16747, B2 => 
                           n16809, ZN => n2581);
   U16978 : OAI22_X1 port map( A1 => n17082, A2 => n16780, B1 => n16748, B2 => 
                           n16809, ZN => n2580);
   U16979 : OAI22_X1 port map( A1 => n17083, A2 => n16780, B1 => n16749, B2 => 
                           n16809, ZN => n2579);
   U16980 : OAI22_X1 port map( A1 => n17159, A2 => n16780, B1 => n16750, B2 => 
                           n16809, ZN => n2578);
   U16981 : OAI22_X1 port map( A1 => n17160, A2 => n16780, B1 => n16751, B2 => 
                           n16807, ZN => n2577);
   U16982 : OAI22_X1 port map( A1 => n17084, A2 => n16780, B1 => n16752, B2 => 
                           n16809, ZN => n2576);
   U16983 : OAI22_X1 port map( A1 => n17085, A2 => n16780, B1 => n16753, B2 => 
                           n16807, ZN => n2575);
   U16984 : OAI22_X1 port map( A1 => n17086, A2 => n16780, B1 => n16754, B2 => 
                           n16809, ZN => n2574);
   U16985 : OAI22_X1 port map( A1 => n17087, A2 => n16780, B1 => n16755, B2 => 
                           n16807, ZN => n2573);
   U16986 : OAI22_X1 port map( A1 => n16954, A2 => n16780, B1 => n16756, B2 => 
                           n16807, ZN => n2572);
   U16987 : OAI22_X1 port map( A1 => n17989, A2 => n16811, B1 => n16757, B2 => 
                           n16809, ZN => n2571);
   U16988 : OAI22_X1 port map( A1 => n17990, A2 => n16780, B1 => n16758, B2 => 
                           n16807, ZN => n2570);
   U16989 : OAI22_X1 port map( A1 => n17991, A2 => n16780, B1 => n16759, B2 => 
                           n16809, ZN => n2569);
   U16990 : OAI22_X1 port map( A1 => n17760, A2 => n16811, B1 => n16760, B2 => 
                           n16807, ZN => n2568);
   U16991 : OAI22_X1 port map( A1 => n17364, A2 => n16811, B1 => n16761, B2 => 
                           n16809, ZN => n2567);
   U16992 : OAI22_X1 port map( A1 => n17365, A2 => n16780, B1 => n16762, B2 => 
                           n16807, ZN => n2566);
   U16993 : OAI22_X1 port map( A1 => n17761, A2 => n16780, B1 => n16763, B2 => 
                           n16809, ZN => n2565);
   U16994 : OAI22_X1 port map( A1 => n17762, A2 => n16811, B1 => n16764, B2 => 
                           n16807, ZN => n2564);
   U16995 : OAI22_X1 port map( A1 => n17763, A2 => n16811, B1 => n16765, B2 => 
                           n16807, ZN => n2563);
   U16996 : OAI22_X1 port map( A1 => n17992, A2 => n16780, B1 => n16766, B2 => 
                           n16807, ZN => n2562);
   U16997 : OAI22_X1 port map( A1 => n17993, A2 => n16780, B1 => n16767, B2 => 
                           n16807, ZN => n2561);
   U16998 : OAI22_X1 port map( A1 => n17994, A2 => n16780, B1 => n16768, B2 => 
                           n16809, ZN => n2560);
   U16999 : OAI22_X1 port map( A1 => n17995, A2 => n16780, B1 => n16769, B2 => 
                           n16807, ZN => n2559);
   U17000 : OAI22_X1 port map( A1 => n17996, A2 => n16811, B1 => n16770, B2 => 
                           n16809, ZN => n2558);
   U17001 : OAI22_X1 port map( A1 => n17366, A2 => n16780, B1 => n16771, B2 => 
                           n16809, ZN => n2557);
   U17002 : OAI22_X1 port map( A1 => n17764, A2 => n16811, B1 => n16772, B2 => 
                           n16809, ZN => n2556);
   U17003 : OAI22_X1 port map( A1 => n17997, A2 => n16780, B1 => n16773, B2 => 
                           n16809, ZN => n2555);
   U17004 : OAI22_X1 port map( A1 => n17998, A2 => n16811, B1 => n16774, B2 => 
                           n16809, ZN => n2554);
   U17005 : OAI22_X1 port map( A1 => n17367, A2 => n16780, B1 => n16775, B2 => 
                           n16809, ZN => n2553);
   U17006 : OAI22_X1 port map( A1 => n17368, A2 => n16811, B1 => n16776, B2 => 
                           n16809, ZN => n2552);
   U17007 : OAI22_X1 port map( A1 => n17369, A2 => n16780, B1 => n16777, B2 => 
                           n16809, ZN => n2551);
   U17008 : OAI22_X1 port map( A1 => n17999, A2 => n16811, B1 => n16778, B2 => 
                           n16809, ZN => n2550);
   U17009 : OAI22_X1 port map( A1 => n18000, A2 => n16780, B1 => n16779, B2 => 
                           n16809, ZN => n2549);
   U17010 : OAI22_X1 port map( A1 => n17765, A2 => n16811, B1 => n16781, B2 => 
                           n16807, ZN => n2548);
   U17011 : OAI22_X1 port map( A1 => n17088, A2 => n16811, B1 => n16782, B2 => 
                           n16807, ZN => n2547);
   U17012 : OAI22_X1 port map( A1 => n16955, A2 => n16780, B1 => n16783, B2 => 
                           n16807, ZN => n2546);
   U17013 : OAI22_X1 port map( A1 => n17161, A2 => n16811, B1 => n16784, B2 => 
                           n16807, ZN => n2545);
   U17014 : OAI22_X1 port map( A1 => n17089, A2 => n16780, B1 => n16785, B2 => 
                           n16807, ZN => n2544);
   U17015 : OAI22_X1 port map( A1 => n17162, A2 => n16811, B1 => n16786, B2 => 
                           n16807, ZN => n2543);
   U17016 : OAI22_X1 port map( A1 => n16956, A2 => n16780, B1 => n16787, B2 => 
                           n16807, ZN => n2542);
   U17017 : OAI22_X1 port map( A1 => n17090, A2 => n16780, B1 => n16788, B2 => 
                           n16807, ZN => n2541);
   U17018 : OAI22_X1 port map( A1 => n17163, A2 => n16780, B1 => n16789, B2 => 
                           n16807, ZN => n2540);
   U17019 : OAI22_X1 port map( A1 => n17091, A2 => n16780, B1 => n16790, B2 => 
                           n16807, ZN => n2539);
   U17020 : OAI22_X1 port map( A1 => n16957, A2 => n16780, B1 => n16791, B2 => 
                           n16807, ZN => n2538);
   U17021 : OAI22_X1 port map( A1 => n17092, A2 => n16780, B1 => n16792, B2 => 
                           n16807, ZN => n2537);
   U17022 : OAI22_X1 port map( A1 => n17164, A2 => n16780, B1 => n16793, B2 => 
                           n16807, ZN => n2536);
   U17023 : OAI22_X1 port map( A1 => n17370, A2 => n16811, B1 => n16794, B2 => 
                           n16807, ZN => n2535);
   U17024 : OAI22_X1 port map( A1 => n17766, A2 => n16811, B1 => n16795, B2 => 
                           n16807, ZN => n2534);
   U17025 : OAI22_X1 port map( A1 => n17371, A2 => n16780, B1 => n16796, B2 => 
                           n16807, ZN => n2533);
   U17026 : OAI22_X1 port map( A1 => n17767, A2 => n16780, B1 => n16797, B2 => 
                           n16807, ZN => n2532);
   U17027 : OAI22_X1 port map( A1 => n17768, A2 => n16811, B1 => n16798, B2 => 
                           n16807, ZN => n2531);
   U17028 : OAI22_X1 port map( A1 => n17372, A2 => n16780, B1 => n16799, B2 => 
                           n16807, ZN => n2530);
   U17029 : OAI22_X1 port map( A1 => n17769, A2 => n16811, B1 => n16800, B2 => 
                           n16807, ZN => n2529);
   U17030 : OAI22_X1 port map( A1 => n17770, A2 => n16780, B1 => n16801, B2 => 
                           n16807, ZN => n2528);
   U17031 : OAI22_X1 port map( A1 => n17771, A2 => n16811, B1 => n16802, B2 => 
                           n16807, ZN => n2527);
   U17032 : OAI22_X1 port map( A1 => n17772, A2 => n16811, B1 => n16803, B2 => 
                           n16807, ZN => n2526);
   U17033 : OAI22_X1 port map( A1 => n18001, A2 => n16780, B1 => n16804, B2 => 
                           n16807, ZN => n2525);
   U17034 : OAI22_X1 port map( A1 => n17773, A2 => n16780, B1 => n16805, B2 => 
                           n16809, ZN => n2524);
   U17035 : OAI22_X1 port map( A1 => n17774, A2 => n16811, B1 => n16806, B2 => 
                           n16807, ZN => n2523);
   U17036 : OAI22_X1 port map( A1 => n17373, A2 => n16780, B1 => n16808, B2 => 
                           n16807, ZN => n2522);
   U17037 : OAI22_X1 port map( A1 => n17775, A2 => n16811, B1 => n16810, B2 => 
                           n16809, ZN => n2521);
   U17038 : OAI22_X1 port map( A1 => n17776, A2 => n16780, B1 => n16812, B2 => 
                           n16807, ZN => n2520);
   U17039 : NAND2_X1 port map( A1 => n16814, A2 => n16813, ZN => n16877);
   U17040 : CLKBUF_X2 port map( A => n16877, Z => n16880);
   U17041 : NAND2_X1 port map( A1 => n13731, A2 => n16880, ZN => n16879);
   U17042 : OAI22_X1 port map( A1 => n18242, A2 => n16879, B1 => n16815, B2 => 
                           n16877, ZN => n2519);
   U17043 : OAI22_X1 port map( A1 => n17093, A2 => n16882, B1 => n16816, B2 => 
                           n16880, ZN => n2518);
   U17044 : OAI22_X1 port map( A1 => n17094, A2 => n16879, B1 => n16817, B2 => 
                           n16877, ZN => n2517);
   U17045 : OAI22_X1 port map( A1 => n16958, A2 => n16882, B1 => n16818, B2 => 
                           n16877, ZN => n2516);
   U17046 : OAI22_X1 port map( A1 => n17165, A2 => n16882, B1 => n16819, B2 => 
                           n16880, ZN => n2515);
   U17047 : OAI22_X1 port map( A1 => n17095, A2 => n16879, B1 => n16820, B2 => 
                           n16877, ZN => n2514);
   U17048 : OAI22_X1 port map( A1 => n16959, A2 => n16882, B1 => n16821, B2 => 
                           n16880, ZN => n2513);
   U17049 : OAI22_X1 port map( A1 => n17166, A2 => n16879, B1 => n16822, B2 => 
                           n16880, ZN => n2512);
   U17050 : OAI22_X1 port map( A1 => n17167, A2 => n16882, B1 => n16823, B2 => 
                           n16880, ZN => n2511);
   U17051 : OAI22_X1 port map( A1 => n17096, A2 => n16879, B1 => n16824, B2 => 
                           n16880, ZN => n2510);
   U17052 : OAI22_X1 port map( A1 => n16960, A2 => n16882, B1 => n16825, B2 => 
                           n16880, ZN => n2509);
   U17053 : OAI22_X1 port map( A1 => n17097, A2 => n16882, B1 => n16826, B2 => 
                           n16877, ZN => n2508);
   U17054 : OAI22_X1 port map( A1 => n17777, A2 => n16879, B1 => n16827, B2 => 
                           n16877, ZN => n2507);
   U17055 : OAI22_X1 port map( A1 => n17778, A2 => n16882, B1 => n16828, B2 => 
                           n16880, ZN => n2506);
   U17056 : OAI22_X1 port map( A1 => n17779, A2 => n16882, B1 => n16829, B2 => 
                           n16877, ZN => n2505);
   U17057 : OAI22_X1 port map( A1 => n18002, A2 => n16879, B1 => n16830, B2 => 
                           n16877, ZN => n2504);
   U17058 : OAI22_X1 port map( A1 => n17374, A2 => n16879, B1 => n16831, B2 => 
                           n16877, ZN => n2503);
   U17059 : OAI22_X1 port map( A1 => n17375, A2 => n16882, B1 => n16832, B2 => 
                           n16880, ZN => n2502);
   U17060 : OAI22_X1 port map( A1 => n17376, A2 => n16882, B1 => n16833, B2 => 
                           n16877, ZN => n2501);
   U17061 : OAI22_X1 port map( A1 => n17377, A2 => n16879, B1 => n16834, B2 => 
                           n16877, ZN => n2500);
   U17062 : OAI22_X1 port map( A1 => n17378, A2 => n16879, B1 => n16835, B2 => 
                           n16880, ZN => n2499);
   U17063 : OAI22_X1 port map( A1 => n17780, A2 => n16882, B1 => n16836, B2 => 
                           n16880, ZN => n2498);
   U17064 : OAI22_X1 port map( A1 => n17379, A2 => n16882, B1 => n16837, B2 => 
                           n16880, ZN => n2497);
   U17065 : OAI22_X1 port map( A1 => n18003, A2 => n16882, B1 => n16838, B2 => 
                           n16877, ZN => n2496);
   U17066 : OAI22_X1 port map( A1 => n17781, A2 => n16882, B1 => n16839, B2 => 
                           n16880, ZN => n2495);
   U17067 : OAI22_X1 port map( A1 => n17782, A2 => n16879, B1 => n16840, B2 => 
                           n16877, ZN => n2494);
   U17068 : OAI22_X1 port map( A1 => n17380, A2 => n16882, B1 => n16841, B2 => 
                           n16877, ZN => n2493);
   U17069 : OAI22_X1 port map( A1 => n17783, A2 => n16879, B1 => n16842, B2 => 
                           n16877, ZN => n2492);
   U17070 : OAI22_X1 port map( A1 => n17784, A2 => n16882, B1 => n16843, B2 => 
                           n16877, ZN => n2491);
   U17071 : OAI22_X1 port map( A1 => n17381, A2 => n16879, B1 => n16844, B2 => 
                           n16877, ZN => n2490);
   U17072 : OAI22_X1 port map( A1 => n17382, A2 => n16882, B1 => n16845, B2 => 
                           n16877, ZN => n2489);
   U17073 : OAI22_X1 port map( A1 => n17383, A2 => n16879, B1 => n16846, B2 => 
                           n16877, ZN => n2488);
   U17074 : OAI22_X1 port map( A1 => n17384, A2 => n16882, B1 => n16847, B2 => 
                           n16877, ZN => n2487);
   U17075 : OAI22_X1 port map( A1 => n17385, A2 => n16879, B1 => n16848, B2 => 
                           n16877, ZN => n2486);
   U17076 : OAI22_X1 port map( A1 => n17785, A2 => n16882, B1 => n16849, B2 => 
                           n16877, ZN => n2485);
   U17077 : OAI22_X1 port map( A1 => n17786, A2 => n16879, B1 => n16850, B2 => 
                           n16880, ZN => n2484);
   U17078 : CLKBUF_X2 port map( A => n16879, Z => n16882);
   U17079 : OAI22_X1 port map( A1 => n17098, A2 => n16882, B1 => n16851, B2 => 
                           n16880, ZN => n2483);
   U17080 : OAI22_X1 port map( A1 => n17099, A2 => n16882, B1 => n16852, B2 => 
                           n16880, ZN => n2482);
   U17081 : OAI22_X1 port map( A1 => n16961, A2 => n16882, B1 => n16853, B2 => 
                           n16880, ZN => n2481);
   U17082 : OAI22_X1 port map( A1 => n17168, A2 => n16882, B1 => n16854, B2 => 
                           n16880, ZN => n2480);
   U17083 : OAI22_X1 port map( A1 => n17100, A2 => n16882, B1 => n16855, B2 => 
                           n16880, ZN => n2479);
   U17084 : OAI22_X1 port map( A1 => n17101, A2 => n16882, B1 => n16856, B2 => 
                           n16880, ZN => n2478);
   U17085 : OAI22_X1 port map( A1 => n17102, A2 => n16882, B1 => n16857, B2 => 
                           n16880, ZN => n2477);
   U17086 : OAI22_X1 port map( A1 => n17103, A2 => n16882, B1 => n16858, B2 => 
                           n16880, ZN => n2476);
   U17087 : OAI22_X1 port map( A1 => n16962, A2 => n16882, B1 => n16859, B2 => 
                           n16880, ZN => n2475);
   U17088 : OAI22_X1 port map( A1 => n17169, A2 => n16882, B1 => n16860, B2 => 
                           n16880, ZN => n2474);
   U17089 : OAI22_X1 port map( A1 => n17104, A2 => n16882, B1 => n16861, B2 => 
                           n16880, ZN => n2473);
   U17090 : OAI22_X1 port map( A1 => n17170, A2 => n16882, B1 => n16862, B2 => 
                           n16880, ZN => n2472);
   U17091 : OAI22_X1 port map( A1 => n17787, A2 => n16879, B1 => n16863, B2 => 
                           n16880, ZN => n2471);
   U17092 : OAI22_X1 port map( A1 => n17386, A2 => n16879, B1 => n16864, B2 => 
                           n16880, ZN => n2470);
   U17093 : OAI22_X1 port map( A1 => n17788, A2 => n16882, B1 => n16865, B2 => 
                           n16880, ZN => n2469);
   U17094 : OAI22_X1 port map( A1 => n18004, A2 => n16882, B1 => n16866, B2 => 
                           n16880, ZN => n2468);
   U17095 : OAI22_X1 port map( A1 => n18005, A2 => n16879, B1 => n16867, B2 => 
                           n16880, ZN => n2467);
   U17096 : OAI22_X1 port map( A1 => n18006, A2 => n16882, B1 => n16868, B2 => 
                           n16880, ZN => n2466);
   U17097 : OAI22_X1 port map( A1 => n18007, A2 => n16879, B1 => n16869, B2 => 
                           n16880, ZN => n2465);
   U17098 : OAI22_X1 port map( A1 => n17789, A2 => n16882, B1 => n16870, B2 => 
                           n16880, ZN => n2464);
   U17099 : OAI22_X1 port map( A1 => n18008, A2 => n16879, B1 => n16871, B2 => 
                           n16880, ZN => n2463);
   U17100 : OAI22_X1 port map( A1 => n17387, A2 => n16879, B1 => n16872, B2 => 
                           n16880, ZN => n2462);
   U17101 : OAI22_X1 port map( A1 => n17790, A2 => n16882, B1 => n16873, B2 => 
                           n16880, ZN => n2461);
   U17102 : OAI22_X1 port map( A1 => n18009, A2 => n16882, B1 => n16874, B2 => 
                           n16877, ZN => n2460);
   U17103 : OAI22_X1 port map( A1 => n18010, A2 => n16879, B1 => n16875, B2 => 
                           n16880, ZN => n2459);
   U17104 : OAI22_X1 port map( A1 => n17791, A2 => n16882, B1 => n16876, B2 => 
                           n16880, ZN => n2458);
   U17105 : OAI22_X1 port map( A1 => n17792, A2 => n16879, B1 => n16878, B2 => 
                           n16877, ZN => n2457);
   U17106 : OAI22_X1 port map( A1 => n17793, A2 => n16882, B1 => n16881, B2 => 
                           n16880, ZN => n2456);

end SYN_A;
