
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_MUX21 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_MUX21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_191 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_191;

architecture SYN_ARCH2 of ND2_191 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_190 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_190;

architecture SYN_ARCH2 of ND2_190 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_189 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_189;

architecture SYN_ARCH2 of ND2_189 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_188 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_188;

architecture SYN_ARCH2 of ND2_188 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_187 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_187;

architecture SYN_ARCH2 of ND2_187 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_186 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_186;

architecture SYN_ARCH2 of ND2_186 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_185 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_185;

architecture SYN_ARCH2 of ND2_185 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_184 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_184;

architecture SYN_ARCH2 of ND2_184 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_183 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_183;

architecture SYN_ARCH2 of ND2_183 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_182 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_182;

architecture SYN_ARCH2 of ND2_182 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_181 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_181;

architecture SYN_ARCH2 of ND2_181 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_180 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_180;

architecture SYN_ARCH2 of ND2_180 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_179 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_179;

architecture SYN_ARCH2 of ND2_179 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_178 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_178;

architecture SYN_ARCH2 of ND2_178 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_177 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_177;

architecture SYN_ARCH2 of ND2_177 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_176 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_176;

architecture SYN_ARCH2 of ND2_176 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_175 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_175;

architecture SYN_ARCH2 of ND2_175 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_174 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_174;

architecture SYN_ARCH2 of ND2_174 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_173 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_173;

architecture SYN_ARCH2 of ND2_173 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_172 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_172;

architecture SYN_ARCH2 of ND2_172 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_171 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_171;

architecture SYN_ARCH2 of ND2_171 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_170 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_170;

architecture SYN_ARCH2 of ND2_170 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_169 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_169;

architecture SYN_ARCH2 of ND2_169 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_168 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_168;

architecture SYN_ARCH2 of ND2_168 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_167 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_167;

architecture SYN_ARCH2 of ND2_167 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_166 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_166;

architecture SYN_ARCH2 of ND2_166 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_165 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_165;

architecture SYN_ARCH2 of ND2_165 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_164 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_164;

architecture SYN_ARCH2 of ND2_164 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_163 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_163;

architecture SYN_ARCH2 of ND2_163 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_162 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_162;

architecture SYN_ARCH2 of ND2_162 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_161 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_161;

architecture SYN_ARCH2 of ND2_161 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_160 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_160;

architecture SYN_ARCH2 of ND2_160 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_159 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_159;

architecture SYN_ARCH2 of ND2_159 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_158 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_158;

architecture SYN_ARCH2 of ND2_158 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_157 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_157;

architecture SYN_ARCH2 of ND2_157 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_156 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_156;

architecture SYN_ARCH2 of ND2_156 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_155 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_155;

architecture SYN_ARCH2 of ND2_155 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_154 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_154;

architecture SYN_ARCH2 of ND2_154 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_153 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_153;

architecture SYN_ARCH2 of ND2_153 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_152 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_152;

architecture SYN_ARCH2 of ND2_152 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_151 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_151;

architecture SYN_ARCH2 of ND2_151 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_150 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_150;

architecture SYN_ARCH2 of ND2_150 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_149 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_149;

architecture SYN_ARCH2 of ND2_149 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_148 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_148;

architecture SYN_ARCH2 of ND2_148 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_147 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_147;

architecture SYN_ARCH2 of ND2_147 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_146 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_146;

architecture SYN_ARCH2 of ND2_146 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_145 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_145;

architecture SYN_ARCH2 of ND2_145 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_144 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_144;

architecture SYN_ARCH2 of ND2_144 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_143 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_143;

architecture SYN_ARCH2 of ND2_143 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_142 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_142;

architecture SYN_ARCH2 of ND2_142 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_141 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_141;

architecture SYN_ARCH2 of ND2_141 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_140 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_140;

architecture SYN_ARCH2 of ND2_140 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_139 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_139;

architecture SYN_ARCH2 of ND2_139 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_138 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_138;

architecture SYN_ARCH2 of ND2_138 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_137 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_137;

architecture SYN_ARCH2 of ND2_137 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_136 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_136;

architecture SYN_ARCH2 of ND2_136 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_135 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_135;

architecture SYN_ARCH2 of ND2_135 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_134 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_134;

architecture SYN_ARCH2 of ND2_134 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_133 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_133;

architecture SYN_ARCH2 of ND2_133 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_132 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_132;

architecture SYN_ARCH2 of ND2_132 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_131 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_131;

architecture SYN_ARCH2 of ND2_131 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_130 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_130;

architecture SYN_ARCH2 of ND2_130 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_129 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_129;

architecture SYN_ARCH2 of ND2_129 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_128 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_128;

architecture SYN_ARCH2 of ND2_128 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_127 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_127;

architecture SYN_ARCH2 of ND2_127 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_126 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_126;

architecture SYN_ARCH2 of ND2_126 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_125 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_125;

architecture SYN_ARCH2 of ND2_125 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_124 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_124;

architecture SYN_ARCH2 of ND2_124 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_123 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_123;

architecture SYN_ARCH2 of ND2_123 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_122 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_122;

architecture SYN_ARCH2 of ND2_122 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_121 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_121;

architecture SYN_ARCH2 of ND2_121 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_120 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_120;

architecture SYN_ARCH2 of ND2_120 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_119 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_119;

architecture SYN_ARCH2 of ND2_119 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_118 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_118;

architecture SYN_ARCH2 of ND2_118 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_117 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_117;

architecture SYN_ARCH2 of ND2_117 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_116 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_116;

architecture SYN_ARCH2 of ND2_116 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_115 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_115;

architecture SYN_ARCH2 of ND2_115 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_114 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_114;

architecture SYN_ARCH2 of ND2_114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_113 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_113;

architecture SYN_ARCH2 of ND2_113 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_112 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_112;

architecture SYN_ARCH2 of ND2_112 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_111 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_111;

architecture SYN_ARCH2 of ND2_111 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_110 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_110;

architecture SYN_ARCH2 of ND2_110 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_109 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_109;

architecture SYN_ARCH2 of ND2_109 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_108 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_108;

architecture SYN_ARCH2 of ND2_108 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_107 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_107;

architecture SYN_ARCH2 of ND2_107 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_106 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_106;

architecture SYN_ARCH2 of ND2_106 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_105 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_105;

architecture SYN_ARCH2 of ND2_105 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_104 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_104;

architecture SYN_ARCH2 of ND2_104 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_103 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_103;

architecture SYN_ARCH2 of ND2_103 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_102 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_102;

architecture SYN_ARCH2 of ND2_102 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_101 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_101;

architecture SYN_ARCH2 of ND2_101 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_100 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_100;

architecture SYN_ARCH2 of ND2_100 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_99 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_99;

architecture SYN_ARCH2 of ND2_99 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_98 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_98;

architecture SYN_ARCH2 of ND2_98 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_97 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_97;

architecture SYN_ARCH2 of ND2_97 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_96 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_96;

architecture SYN_ARCH2 of ND2_96 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_95 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_95;

architecture SYN_ARCH2 of ND2_95 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_94 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_94;

architecture SYN_ARCH2 of ND2_94 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_93 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_93;

architecture SYN_ARCH2 of ND2_93 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_92 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_92;

architecture SYN_ARCH2 of ND2_92 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_91 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_91;

architecture SYN_ARCH2 of ND2_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_90 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_90;

architecture SYN_ARCH2 of ND2_90 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_89 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_89;

architecture SYN_ARCH2 of ND2_89 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_88 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_88;

architecture SYN_ARCH2 of ND2_88 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_87 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_87;

architecture SYN_ARCH2 of ND2_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_86 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_86;

architecture SYN_ARCH2 of ND2_86 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_85 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_85;

architecture SYN_ARCH2 of ND2_85 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_84 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_84;

architecture SYN_ARCH2 of ND2_84 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_83 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_83;

architecture SYN_ARCH2 of ND2_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_82 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_82;

architecture SYN_ARCH2 of ND2_82 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_81 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_81;

architecture SYN_ARCH2 of ND2_81 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_80 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_80;

architecture SYN_ARCH2 of ND2_80 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_79 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_79;

architecture SYN_ARCH2 of ND2_79 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_78 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_78;

architecture SYN_ARCH2 of ND2_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_77 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_77;

architecture SYN_ARCH2 of ND2_77 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_76 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_76;

architecture SYN_ARCH2 of ND2_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_75 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_75;

architecture SYN_ARCH2 of ND2_75 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_74 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_74;

architecture SYN_ARCH2 of ND2_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_73 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_73;

architecture SYN_ARCH2 of ND2_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_72 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_72;

architecture SYN_ARCH2 of ND2_72 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_71 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_71;

architecture SYN_ARCH2 of ND2_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_70 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_70;

architecture SYN_ARCH2 of ND2_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_69 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_69;

architecture SYN_ARCH2 of ND2_69 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_68 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_68;

architecture SYN_ARCH2 of ND2_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_67 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_67;

architecture SYN_ARCH2 of ND2_67 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_66 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_66;

architecture SYN_ARCH2 of ND2_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_65 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_65;

architecture SYN_ARCH2 of ND2_65 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_64 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_64;

architecture SYN_ARCH2 of ND2_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_63;

architecture SYN_ARCH2 of ND2_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_62;

architecture SYN_ARCH2 of ND2_62 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_61;

architecture SYN_ARCH2 of ND2_61 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_60;

architecture SYN_ARCH2 of ND2_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_59;

architecture SYN_ARCH2 of ND2_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_58;

architecture SYN_ARCH2 of ND2_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_57;

architecture SYN_ARCH2 of ND2_57 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_56;

architecture SYN_ARCH2 of ND2_56 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_55;

architecture SYN_ARCH2 of ND2_55 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_54;

architecture SYN_ARCH2 of ND2_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_53;

architecture SYN_ARCH2 of ND2_53 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_52;

architecture SYN_ARCH2 of ND2_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_51;

architecture SYN_ARCH2 of ND2_51 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_50;

architecture SYN_ARCH2 of ND2_50 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_49;

architecture SYN_ARCH2 of ND2_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_48;

architecture SYN_ARCH2 of ND2_48 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_47;

architecture SYN_ARCH2 of ND2_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_46;

architecture SYN_ARCH2 of ND2_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_45;

architecture SYN_ARCH2 of ND2_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_44;

architecture SYN_ARCH2 of ND2_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_43;

architecture SYN_ARCH2 of ND2_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_42;

architecture SYN_ARCH2 of ND2_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_41;

architecture SYN_ARCH2 of ND2_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_40;

architecture SYN_ARCH2 of ND2_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_39;

architecture SYN_ARCH2 of ND2_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_38;

architecture SYN_ARCH2 of ND2_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_37;

architecture SYN_ARCH2 of ND2_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_36;

architecture SYN_ARCH2 of ND2_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_35;

architecture SYN_ARCH2 of ND2_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_34;

architecture SYN_ARCH2 of ND2_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_33;

architecture SYN_ARCH2 of ND2_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_32;

architecture SYN_ARCH2 of ND2_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_31;

architecture SYN_ARCH2 of ND2_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_30;

architecture SYN_ARCH2 of ND2_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_29;

architecture SYN_ARCH2 of ND2_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_28;

architecture SYN_ARCH2 of ND2_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_27;

architecture SYN_ARCH2 of ND2_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_26;

architecture SYN_ARCH2 of ND2_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_25;

architecture SYN_ARCH2 of ND2_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_24;

architecture SYN_ARCH2 of ND2_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_23;

architecture SYN_ARCH2 of ND2_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_22;

architecture SYN_ARCH2 of ND2_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_21;

architecture SYN_ARCH2 of ND2_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_20;

architecture SYN_ARCH2 of ND2_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_19;

architecture SYN_ARCH2 of ND2_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_18;

architecture SYN_ARCH2 of ND2_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_17;

architecture SYN_ARCH2 of ND2_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_16;

architecture SYN_ARCH2 of ND2_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_15;

architecture SYN_ARCH2 of ND2_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_14;

architecture SYN_ARCH2 of ND2_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_13;

architecture SYN_ARCH2 of ND2_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_12;

architecture SYN_ARCH2 of ND2_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_11;

architecture SYN_ARCH2 of ND2_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_10;

architecture SYN_ARCH2 of ND2_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_9;

architecture SYN_ARCH2 of ND2_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_8;

architecture SYN_ARCH2 of ND2_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_7;

architecture SYN_ARCH2 of ND2_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_6;

architecture SYN_ARCH2 of ND2_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_5;

architecture SYN_ARCH2 of ND2_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_4;

architecture SYN_ARCH2 of ND2_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_3;

architecture SYN_ARCH2 of ND2_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_2;

architecture SYN_ARCH2 of ND2_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_1;

architecture SYN_ARCH2 of ND2_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity ND2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_0;

architecture SYN_ARCH2 of ND2_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity IV is

   port( A : in std_logic;  Y : out std_logic);

end IV;

architecture SYN_BEHAVIORAL of IV is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21.all;

entity MUX21 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21;

architecture SYN_STRUCTURAL of MUX21 is

   component ND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_64
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_65
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_66
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_67
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_68
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_69
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_70
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_71
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_72
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_73
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_74
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_75
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_76
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_77
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_78
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_79
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_80
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_81
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_82
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_83
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_84
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_85
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_86
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_87
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_88
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_89
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_90
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_91
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_92
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_93
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_94
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_95
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_96
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_97
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_98
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_99
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_100
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_101
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_102
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_103
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_104
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_105
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_106
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_107
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_108
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_109
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_110
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_111
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_112
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_113
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_114
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_115
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_116
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_117
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_118
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_119
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_120
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_121
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_122
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_123
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_124
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_125
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_126
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_127
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_128
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_129
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_130
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_131
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_132
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_133
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_134
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_135
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_136
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_137
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_138
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_139
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_140
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_141
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_142
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_143
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_144
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_145
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_146
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_147
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_148
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_149
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_150
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_151
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_152
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_153
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_154
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_155
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_156
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_157
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_158
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_159
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_160
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_161
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_162
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_163
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_164
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_165
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_166
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_167
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_168
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_169
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_170
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_171
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_172
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_173
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_174
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_175
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_176
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_177
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_178
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_179
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_180
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_181
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_182
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_183
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_184
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_185
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_186
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_187
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_188
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_189
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_190
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_191
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal A_S_63_port, A_S_62_port, A_S_61_port, A_S_60_port, A_S_59_port, 
      A_S_58_port, A_S_57_port, A_S_56_port, A_S_55_port, A_S_54_port, 
      A_S_53_port, A_S_52_port, A_S_51_port, A_S_50_port, A_S_49_port, 
      A_S_48_port, A_S_47_port, A_S_46_port, A_S_45_port, A_S_44_port, 
      A_S_43_port, A_S_42_port, A_S_41_port, A_S_40_port, A_S_39_port, 
      A_S_38_port, A_S_37_port, A_S_36_port, A_S_35_port, A_S_34_port, 
      A_S_33_port, A_S_32_port, A_S_31_port, A_S_30_port, A_S_29_port, 
      A_S_28_port, A_S_27_port, A_S_26_port, A_S_25_port, A_S_24_port, 
      A_S_23_port, A_S_22_port, A_S_21_port, A_S_20_port, A_S_19_port, 
      A_S_18_port, A_S_17_port, A_S_16_port, A_S_15_port, A_S_14_port, 
      A_S_13_port, A_S_12_port, A_S_11_port, A_S_10_port, A_S_9_port, 
      A_S_8_port, A_S_7_port, A_S_6_port, A_S_5_port, A_S_4_port, A_S_3_port, 
      A_S_2_port, A_S_1_port, A_S_0_port, B_S_63_port, B_S_62_port, B_S_61_port
      , B_S_60_port, B_S_59_port, B_S_58_port, B_S_57_port, B_S_56_port, 
      B_S_55_port, B_S_54_port, B_S_53_port, B_S_52_port, B_S_51_port, 
      B_S_50_port, B_S_49_port, B_S_48_port, B_S_47_port, B_S_46_port, 
      B_S_45_port, B_S_44_port, B_S_43_port, B_S_42_port, B_S_41_port, 
      B_S_40_port, B_S_39_port, B_S_38_port, B_S_37_port, B_S_36_port, 
      B_S_35_port, B_S_34_port, B_S_33_port, B_S_32_port, B_S_31_port, 
      B_S_30_port, B_S_29_port, B_S_28_port, B_S_27_port, B_S_26_port, 
      B_S_25_port, B_S_24_port, B_S_23_port, B_S_22_port, B_S_21_port, 
      B_S_20_port, B_S_19_port, B_S_18_port, B_S_17_port, B_S_16_port, 
      B_S_15_port, B_S_14_port, B_S_13_port, B_S_12_port, B_S_11_port, 
      B_S_10_port, B_S_9_port, B_S_8_port, B_S_7_port, B_S_6_port, B_S_5_port, 
      B_S_4_port, B_S_3_port, B_S_2_port, B_S_1_port, B_S_0_port, n_1000 : 
      std_logic;

begin
   
   INV : IV port map( A => SEL, Y => n_1000);
   r1_0 : ND2_0 port map( A => A(0), B => SEL, Y => A_S_0_port);
   r1_1 : ND2_191 port map( A => A(1), B => SEL, Y => A_S_1_port);
   r1_2 : ND2_190 port map( A => A(2), B => SEL, Y => A_S_2_port);
   r1_3 : ND2_189 port map( A => A(3), B => SEL, Y => A_S_3_port);
   r1_4 : ND2_188 port map( A => A(4), B => SEL, Y => A_S_4_port);
   r1_5 : ND2_187 port map( A => A(5), B => SEL, Y => A_S_5_port);
   r1_6 : ND2_186 port map( A => A(6), B => SEL, Y => A_S_6_port);
   r1_7 : ND2_185 port map( A => A(7), B => SEL, Y => A_S_7_port);
   r1_8 : ND2_184 port map( A => A(8), B => SEL, Y => A_S_8_port);
   r1_9 : ND2_183 port map( A => A(9), B => SEL, Y => A_S_9_port);
   r1_10 : ND2_182 port map( A => A(10), B => SEL, Y => A_S_10_port);
   r1_11 : ND2_181 port map( A => A(11), B => SEL, Y => A_S_11_port);
   r1_12 : ND2_180 port map( A => A(12), B => SEL, Y => A_S_12_port);
   r1_13 : ND2_179 port map( A => A(13), B => SEL, Y => A_S_13_port);
   r1_14 : ND2_178 port map( A => A(14), B => SEL, Y => A_S_14_port);
   r1_15 : ND2_177 port map( A => A(15), B => SEL, Y => A_S_15_port);
   r1_16 : ND2_176 port map( A => A(16), B => SEL, Y => A_S_16_port);
   r1_17 : ND2_175 port map( A => A(17), B => SEL, Y => A_S_17_port);
   r1_18 : ND2_174 port map( A => A(18), B => SEL, Y => A_S_18_port);
   r1_19 : ND2_173 port map( A => A(19), B => SEL, Y => A_S_19_port);
   r1_20 : ND2_172 port map( A => A(20), B => SEL, Y => A_S_20_port);
   r1_21 : ND2_171 port map( A => A(21), B => SEL, Y => A_S_21_port);
   r1_22 : ND2_170 port map( A => A(22), B => SEL, Y => A_S_22_port);
   r1_23 : ND2_169 port map( A => A(23), B => SEL, Y => A_S_23_port);
   r1_24 : ND2_168 port map( A => A(24), B => SEL, Y => A_S_24_port);
   r1_25 : ND2_167 port map( A => A(25), B => SEL, Y => A_S_25_port);
   r1_26 : ND2_166 port map( A => A(26), B => SEL, Y => A_S_26_port);
   r1_27 : ND2_165 port map( A => A(27), B => SEL, Y => A_S_27_port);
   r1_28 : ND2_164 port map( A => A(28), B => SEL, Y => A_S_28_port);
   r1_29 : ND2_163 port map( A => A(29), B => SEL, Y => A_S_29_port);
   r1_30 : ND2_162 port map( A => A(30), B => SEL, Y => A_S_30_port);
   r1_31 : ND2_161 port map( A => A(31), B => SEL, Y => A_S_31_port);
   r1_32 : ND2_160 port map( A => A(32), B => SEL, Y => A_S_32_port);
   r1_33 : ND2_159 port map( A => A(33), B => SEL, Y => A_S_33_port);
   r1_34 : ND2_158 port map( A => A(34), B => SEL, Y => A_S_34_port);
   r1_35 : ND2_157 port map( A => A(35), B => SEL, Y => A_S_35_port);
   r1_36 : ND2_156 port map( A => A(36), B => SEL, Y => A_S_36_port);
   r1_37 : ND2_155 port map( A => A(37), B => SEL, Y => A_S_37_port);
   r1_38 : ND2_154 port map( A => A(38), B => SEL, Y => A_S_38_port);
   r1_39 : ND2_153 port map( A => A(39), B => SEL, Y => A_S_39_port);
   r1_40 : ND2_152 port map( A => A(40), B => SEL, Y => A_S_40_port);
   r1_41 : ND2_151 port map( A => A(41), B => SEL, Y => A_S_41_port);
   r1_42 : ND2_150 port map( A => A(42), B => SEL, Y => A_S_42_port);
   r1_43 : ND2_149 port map( A => A(43), B => SEL, Y => A_S_43_port);
   r1_44 : ND2_148 port map( A => A(44), B => SEL, Y => A_S_44_port);
   r1_45 : ND2_147 port map( A => A(45), B => SEL, Y => A_S_45_port);
   r1_46 : ND2_146 port map( A => A(46), B => SEL, Y => A_S_46_port);
   r1_47 : ND2_145 port map( A => A(47), B => SEL, Y => A_S_47_port);
   r1_48 : ND2_144 port map( A => A(48), B => SEL, Y => A_S_48_port);
   r1_49 : ND2_143 port map( A => A(49), B => SEL, Y => A_S_49_port);
   r1_50 : ND2_142 port map( A => A(50), B => SEL, Y => A_S_50_port);
   r1_51 : ND2_141 port map( A => A(51), B => SEL, Y => A_S_51_port);
   r1_52 : ND2_140 port map( A => A(52), B => SEL, Y => A_S_52_port);
   r1_53 : ND2_139 port map( A => A(53), B => SEL, Y => A_S_53_port);
   r1_54 : ND2_138 port map( A => A(54), B => SEL, Y => A_S_54_port);
   r1_55 : ND2_137 port map( A => A(55), B => SEL, Y => A_S_55_port);
   r1_56 : ND2_136 port map( A => A(56), B => SEL, Y => A_S_56_port);
   r1_57 : ND2_135 port map( A => A(57), B => SEL, Y => A_S_57_port);
   r1_58 : ND2_134 port map( A => A(58), B => SEL, Y => A_S_58_port);
   r1_59 : ND2_133 port map( A => A(59), B => SEL, Y => A_S_59_port);
   r1_60 : ND2_132 port map( A => A(60), B => SEL, Y => A_S_60_port);
   r1_61 : ND2_131 port map( A => A(61), B => SEL, Y => A_S_61_port);
   r1_62 : ND2_130 port map( A => A(62), B => SEL, Y => A_S_62_port);
   r1_63 : ND2_129 port map( A => A(63), B => SEL, Y => A_S_63_port);
   r2_0 : ND2_128 port map( A => B(0), B => SEL, Y => B_S_0_port);
   r2_1 : ND2_127 port map( A => B(1), B => SEL, Y => B_S_1_port);
   r2_2 : ND2_126 port map( A => B(2), B => SEL, Y => B_S_2_port);
   r2_3 : ND2_125 port map( A => B(3), B => SEL, Y => B_S_3_port);
   r2_4 : ND2_124 port map( A => B(4), B => SEL, Y => B_S_4_port);
   r2_5 : ND2_123 port map( A => B(5), B => SEL, Y => B_S_5_port);
   r2_6 : ND2_122 port map( A => B(6), B => SEL, Y => B_S_6_port);
   r2_7 : ND2_121 port map( A => B(7), B => SEL, Y => B_S_7_port);
   r2_8 : ND2_120 port map( A => B(8), B => SEL, Y => B_S_8_port);
   r2_9 : ND2_119 port map( A => B(9), B => SEL, Y => B_S_9_port);
   r2_10 : ND2_118 port map( A => B(10), B => SEL, Y => B_S_10_port);
   r2_11 : ND2_117 port map( A => B(11), B => SEL, Y => B_S_11_port);
   r2_12 : ND2_116 port map( A => B(12), B => SEL, Y => B_S_12_port);
   r2_13 : ND2_115 port map( A => B(13), B => SEL, Y => B_S_13_port);
   r2_14 : ND2_114 port map( A => B(14), B => SEL, Y => B_S_14_port);
   r2_15 : ND2_113 port map( A => B(15), B => SEL, Y => B_S_15_port);
   r2_16 : ND2_112 port map( A => B(16), B => SEL, Y => B_S_16_port);
   r2_17 : ND2_111 port map( A => B(17), B => SEL, Y => B_S_17_port);
   r2_18 : ND2_110 port map( A => B(18), B => SEL, Y => B_S_18_port);
   r2_19 : ND2_109 port map( A => B(19), B => SEL, Y => B_S_19_port);
   r2_20 : ND2_108 port map( A => B(20), B => SEL, Y => B_S_20_port);
   r2_21 : ND2_107 port map( A => B(21), B => SEL, Y => B_S_21_port);
   r2_22 : ND2_106 port map( A => B(22), B => SEL, Y => B_S_22_port);
   r2_23 : ND2_105 port map( A => B(23), B => SEL, Y => B_S_23_port);
   r2_24 : ND2_104 port map( A => B(24), B => SEL, Y => B_S_24_port);
   r2_25 : ND2_103 port map( A => B(25), B => SEL, Y => B_S_25_port);
   r2_26 : ND2_102 port map( A => B(26), B => SEL, Y => B_S_26_port);
   r2_27 : ND2_101 port map( A => B(27), B => SEL, Y => B_S_27_port);
   r2_28 : ND2_100 port map( A => B(28), B => SEL, Y => B_S_28_port);
   r2_29 : ND2_99 port map( A => B(29), B => SEL, Y => B_S_29_port);
   r2_30 : ND2_98 port map( A => B(30), B => SEL, Y => B_S_30_port);
   r2_31 : ND2_97 port map( A => B(31), B => SEL, Y => B_S_31_port);
   r2_32 : ND2_96 port map( A => B(32), B => SEL, Y => B_S_32_port);
   r2_33 : ND2_95 port map( A => B(33), B => SEL, Y => B_S_33_port);
   r2_34 : ND2_94 port map( A => B(34), B => SEL, Y => B_S_34_port);
   r2_35 : ND2_93 port map( A => B(35), B => SEL, Y => B_S_35_port);
   r2_36 : ND2_92 port map( A => B(36), B => SEL, Y => B_S_36_port);
   r2_37 : ND2_91 port map( A => B(37), B => SEL, Y => B_S_37_port);
   r2_38 : ND2_90 port map( A => B(38), B => SEL, Y => B_S_38_port);
   r2_39 : ND2_89 port map( A => B(39), B => SEL, Y => B_S_39_port);
   r2_40 : ND2_88 port map( A => B(40), B => SEL, Y => B_S_40_port);
   r2_41 : ND2_87 port map( A => B(41), B => SEL, Y => B_S_41_port);
   r2_42 : ND2_86 port map( A => B(42), B => SEL, Y => B_S_42_port);
   r2_43 : ND2_85 port map( A => B(43), B => SEL, Y => B_S_43_port);
   r2_44 : ND2_84 port map( A => B(44), B => SEL, Y => B_S_44_port);
   r2_45 : ND2_83 port map( A => B(45), B => SEL, Y => B_S_45_port);
   r2_46 : ND2_82 port map( A => B(46), B => SEL, Y => B_S_46_port);
   r2_47 : ND2_81 port map( A => B(47), B => SEL, Y => B_S_47_port);
   r2_48 : ND2_80 port map( A => B(48), B => SEL, Y => B_S_48_port);
   r2_49 : ND2_79 port map( A => B(49), B => SEL, Y => B_S_49_port);
   r2_50 : ND2_78 port map( A => B(50), B => SEL, Y => B_S_50_port);
   r2_51 : ND2_77 port map( A => B(51), B => SEL, Y => B_S_51_port);
   r2_52 : ND2_76 port map( A => B(52), B => SEL, Y => B_S_52_port);
   r2_53 : ND2_75 port map( A => B(53), B => SEL, Y => B_S_53_port);
   r2_54 : ND2_74 port map( A => B(54), B => SEL, Y => B_S_54_port);
   r2_55 : ND2_73 port map( A => B(55), B => SEL, Y => B_S_55_port);
   r2_56 : ND2_72 port map( A => B(56), B => SEL, Y => B_S_56_port);
   r2_57 : ND2_71 port map( A => B(57), B => SEL, Y => B_S_57_port);
   r2_58 : ND2_70 port map( A => B(58), B => SEL, Y => B_S_58_port);
   r2_59 : ND2_69 port map( A => B(59), B => SEL, Y => B_S_59_port);
   r2_60 : ND2_68 port map( A => B(60), B => SEL, Y => B_S_60_port);
   r2_61 : ND2_67 port map( A => B(61), B => SEL, Y => B_S_61_port);
   r2_62 : ND2_66 port map( A => B(62), B => SEL, Y => B_S_62_port);
   r2_63 : ND2_65 port map( A => B(63), B => SEL, Y => B_S_63_port);
   r4_0 : ND2_64 port map( A => A_S_0_port, B => B_S_0_port, Y => Y(0));
   r4_1 : ND2_63 port map( A => A_S_1_port, B => B_S_1_port, Y => Y(1));
   r4_2 : ND2_62 port map( A => A_S_2_port, B => B_S_2_port, Y => Y(2));
   r4_3 : ND2_61 port map( A => A_S_3_port, B => B_S_3_port, Y => Y(3));
   r4_4 : ND2_60 port map( A => A_S_4_port, B => B_S_4_port, Y => Y(4));
   r4_5 : ND2_59 port map( A => A_S_5_port, B => B_S_5_port, Y => Y(5));
   r4_6 : ND2_58 port map( A => A_S_6_port, B => B_S_6_port, Y => Y(6));
   r4_7 : ND2_57 port map( A => A_S_7_port, B => B_S_7_port, Y => Y(7));
   r4_8 : ND2_56 port map( A => A_S_8_port, B => B_S_8_port, Y => Y(8));
   r4_9 : ND2_55 port map( A => A_S_9_port, B => B_S_9_port, Y => Y(9));
   r4_10 : ND2_54 port map( A => A_S_10_port, B => B_S_10_port, Y => Y(10));
   r4_11 : ND2_53 port map( A => A_S_11_port, B => B_S_11_port, Y => Y(11));
   r4_12 : ND2_52 port map( A => A_S_12_port, B => B_S_12_port, Y => Y(12));
   r4_13 : ND2_51 port map( A => A_S_13_port, B => B_S_13_port, Y => Y(13));
   r4_14 : ND2_50 port map( A => A_S_14_port, B => B_S_14_port, Y => Y(14));
   r4_15 : ND2_49 port map( A => A_S_15_port, B => B_S_15_port, Y => Y(15));
   r4_16 : ND2_48 port map( A => A_S_16_port, B => B_S_16_port, Y => Y(16));
   r4_17 : ND2_47 port map( A => A_S_17_port, B => B_S_17_port, Y => Y(17));
   r4_18 : ND2_46 port map( A => A_S_18_port, B => B_S_18_port, Y => Y(18));
   r4_19 : ND2_45 port map( A => A_S_19_port, B => B_S_19_port, Y => Y(19));
   r4_20 : ND2_44 port map( A => A_S_20_port, B => B_S_20_port, Y => Y(20));
   r4_21 : ND2_43 port map( A => A_S_21_port, B => B_S_21_port, Y => Y(21));
   r4_22 : ND2_42 port map( A => A_S_22_port, B => B_S_22_port, Y => Y(22));
   r4_23 : ND2_41 port map( A => A_S_23_port, B => B_S_23_port, Y => Y(23));
   r4_24 : ND2_40 port map( A => A_S_24_port, B => B_S_24_port, Y => Y(24));
   r4_25 : ND2_39 port map( A => A_S_25_port, B => B_S_25_port, Y => Y(25));
   r4_26 : ND2_38 port map( A => A_S_26_port, B => B_S_26_port, Y => Y(26));
   r4_27 : ND2_37 port map( A => A_S_27_port, B => B_S_27_port, Y => Y(27));
   r4_28 : ND2_36 port map( A => A_S_28_port, B => B_S_28_port, Y => Y(28));
   r4_29 : ND2_35 port map( A => A_S_29_port, B => B_S_29_port, Y => Y(29));
   r4_30 : ND2_34 port map( A => A_S_30_port, B => B_S_30_port, Y => Y(30));
   r4_31 : ND2_33 port map( A => A_S_31_port, B => B_S_31_port, Y => Y(31));
   r4_32 : ND2_32 port map( A => A_S_32_port, B => B_S_32_port, Y => Y(32));
   r4_33 : ND2_31 port map( A => A_S_33_port, B => B_S_33_port, Y => Y(33));
   r4_34 : ND2_30 port map( A => A_S_34_port, B => B_S_34_port, Y => Y(34));
   r4_35 : ND2_29 port map( A => A_S_35_port, B => B_S_35_port, Y => Y(35));
   r4_36 : ND2_28 port map( A => A_S_36_port, B => B_S_36_port, Y => Y(36));
   r4_37 : ND2_27 port map( A => A_S_37_port, B => B_S_37_port, Y => Y(37));
   r4_38 : ND2_26 port map( A => A_S_38_port, B => B_S_38_port, Y => Y(38));
   r4_39 : ND2_25 port map( A => A_S_39_port, B => B_S_39_port, Y => Y(39));
   r4_40 : ND2_24 port map( A => A_S_40_port, B => B_S_40_port, Y => Y(40));
   r4_41 : ND2_23 port map( A => A_S_41_port, B => B_S_41_port, Y => Y(41));
   r4_42 : ND2_22 port map( A => A_S_42_port, B => B_S_42_port, Y => Y(42));
   r4_43 : ND2_21 port map( A => A_S_43_port, B => B_S_43_port, Y => Y(43));
   r4_44 : ND2_20 port map( A => A_S_44_port, B => B_S_44_port, Y => Y(44));
   r4_45 : ND2_19 port map( A => A_S_45_port, B => B_S_45_port, Y => Y(45));
   r4_46 : ND2_18 port map( A => A_S_46_port, B => B_S_46_port, Y => Y(46));
   r4_47 : ND2_17 port map( A => A_S_47_port, B => B_S_47_port, Y => Y(47));
   r4_48 : ND2_16 port map( A => A_S_48_port, B => B_S_48_port, Y => Y(48));
   r4_49 : ND2_15 port map( A => A_S_49_port, B => B_S_49_port, Y => Y(49));
   r4_50 : ND2_14 port map( A => A_S_50_port, B => B_S_50_port, Y => Y(50));
   r4_51 : ND2_13 port map( A => A_S_51_port, B => B_S_51_port, Y => Y(51));
   r4_52 : ND2_12 port map( A => A_S_52_port, B => B_S_52_port, Y => Y(52));
   r4_53 : ND2_11 port map( A => A_S_53_port, B => B_S_53_port, Y => Y(53));
   r4_54 : ND2_10 port map( A => A_S_54_port, B => B_S_54_port, Y => Y(54));
   r4_55 : ND2_9 port map( A => A_S_55_port, B => B_S_55_port, Y => Y(55));
   r4_56 : ND2_8 port map( A => A_S_56_port, B => B_S_56_port, Y => Y(56));
   r4_57 : ND2_7 port map( A => A_S_57_port, B => B_S_57_port, Y => Y(57));
   r4_58 : ND2_6 port map( A => A_S_58_port, B => B_S_58_port, Y => Y(58));
   r4_59 : ND2_5 port map( A => A_S_59_port, B => B_S_59_port, Y => Y(59));
   r4_60 : ND2_4 port map( A => A_S_60_port, B => B_S_60_port, Y => Y(60));
   r4_61 : ND2_3 port map( A => A_S_61_port, B => B_S_61_port, Y => Y(61));
   r4_62 : ND2_2 port map( A => A_S_62_port, B => B_S_62_port, Y => Y(62));
   r4_63 : ND2_1 port map( A => A_S_63_port, B => B_S_63_port, Y => Y(63));

end SYN_STRUCTURAL;
